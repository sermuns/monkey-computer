LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY pMem IS
    PORT (
        clk : IN STD_LOGIC;
        cpu_address : IN unsigned(11 DOWNTO 0);
        cpu_data_out : OUT STD_LOGIC_VECTOR(23 DOWNTO 0);
        cpu_data_in : IN unsigned(23 DOWNTO 0);
        cpu_we : IN STD_LOGIC;
        video_address : IN unsigned(6 DOWNTO 0);
        video_data : OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
    );
END pMem;

ARCHITECTURE func OF pMem IS

    TYPE p_mem_type IS ARRAY(0 TO 4095) OF STD_LOGIC_VECTOR(23 DOWNTO 0);

    CONSTANT PROGRAM : INTEGER := 0;
    CONSTANT VMEM : INTEGER := 1500;
    CONSTANT PATH : INTEGER := 1600;
    CONSTANT HEAP : INTEGER := 3000;

    -- 00000_000_00_00_000000000000
    -- OP    GRx M  *  ADR 
    -- 5     3   2  2  12  
    SIGNAL p_mem : p_mem_type := (
        -- PROGRAM
        PROGRAM + 0 => b"01010_000_00_00_000000000000", -- BRA :
        PROGRAM + 1 => b"01010_000_00_00_000000000000", -- BRA :
        PROGRAM + 2 => b"11111_---_--_--_------------", -- HALT : 
        -- VMEM
        VMEM + 0 => b"000000000000000000000000", -- 0 : 
        VMEM + 1 => b"000000000000000000000000", -- 0 : 
        VMEM + 2 => b"000000000000000000000000", -- 0 : 
        VMEM + 3 => b"000000000000000000000000", -- 0 : 
        VMEM + 4 => b"000000000000000000000000", -- 0 : 
        VMEM + 5 => b"000000000000000000000000", -- 0 : 
        VMEM + 6 => b"000000000000000000000010", -- 0 : 
        VMEM + 7 => b"000000000000000000000000", -- 0 : 
        VMEM + 8 => b"000000000000000000000000", -- 0 : 
        VMEM + 9 => b"000000000000000000000101", -- 0 : 
        VMEM + 10 => b"000000000000000000000000", -- 0 : 
        VMEM + 11 => b"000000000000000000011001", -- 25 : 
        VMEM + 12 => b"000000000000000000011001", -- 25 : 
        VMEM + 13 => b"000000000000000000011001", -- 25 : 
        VMEM + 14 => b"000000000000000000011001", -- 25 : 
        VMEM + 15 => b"000000000000000000011001", -- 25 : 
        VMEM + 16 => b"000000000000000000011001", -- 25 : 
        VMEM + 17 => b"000000000000000000011001", -- 25 : 
        VMEM + 18 => b"000000000000000000011001", -- 25 : 
        VMEM + 19 => b"000000000000000000000000", -- 0 : 
        VMEM + 20 => b"000000000000000000000000", -- 0 : 
        VMEM + 21 => b"000000000000000000011001", -- 25 : 
        VMEM + 22 => b"000000000000000000000000", -- 0 : 
        VMEM + 23 => b"000000000000000000000000", -- 0 : 
        VMEM + 24 => b"000000000000000000000000", -- 0 : 
        VMEM + 25 => b"000000000000000000000000", -- 0 : 
        VMEM + 26 => b"000000000000000000000000", -- 0 : 
        VMEM + 27 => b"000000000000000000000000", -- 0 : 
        VMEM + 28 => b"000000000000000000011001", -- 25 : 
        VMEM + 29 => b"000000000000000000000000", -- 0 : 
        VMEM + 30 => b"000000000000000000000000", -- 0 : 
        VMEM + 31 => b"000000000000000000011001", -- 25 : 
        VMEM + 32 => b"000000000000000000000000", -- 0 : 
        VMEM + 33 => b"000000000000000000011001", -- 25 : 
        VMEM + 34 => b"000000000000000000011001", -- 25 : 
        VMEM + 35 => b"000000000000000000011001", -- 25 : 
        VMEM + 36 => b"000000000000000000011001", -- 25 : 
        VMEM + 37 => b"000000000000000000011001", -- 25 : 
        VMEM + 38 => b"000000000000000000011001", -- 25 : 
        VMEM + 39 => b"000000000000000000000000", -- 0 : 
        VMEM + 40 => b"000000000000000000011001", -- 25 : 
        VMEM + 41 => b"000000000000000000011001", -- 25 : 
        VMEM + 42 => b"000000000000000000000000", -- 0 : 
        VMEM + 43 => b"000000000000000000011001", -- 25 : 
        VMEM + 44 => b"000000000000000000000000", -- 0 : 
        VMEM + 45 => b"000000000000000000000000", -- 0 : 
        VMEM + 46 => b"000000000000000000000000", -- 0 : 
        VMEM + 47 => b"000000000000000000000000", -- 0 : 
        VMEM + 48 => b"000000000000000000000000", -- 0 : 
        VMEM + 49 => b"000000000000000000000000", -- 0 : 
        VMEM + 50 => b"000000000000000000000000", -- 0 : 
        VMEM + 51 => b"000000000000000000000000", -- 0 : 
        VMEM + 52 => b"000000000000000000000000", -- 0 : 
        VMEM + 53 => b"000000000000000000011001", -- 25 : 
        VMEM + 54 => b"000000000000000000000000", -- 0 : 
        VMEM + 55 => b"000000000000000000011001", -- 25 : 
        VMEM + 56 => b"000000000000000000011001", -- 25 : 
        VMEM + 57 => b"000000000000000000011001", -- 25 : 
        VMEM + 58 => b"000000000000000000000000", -- 0 : 
        VMEM + 59 => b"000000000000000000000000", -- 0 : 
        VMEM + 60 => b"000000000000000000000000", -- 0 : 
        VMEM + 61 => b"000000000000000000011001", -- 25 : 
        VMEM + 62 => b"000000000000000000011001", -- 25 : 
        VMEM + 63 => b"000000000000000000011001", -- 25 : 
        VMEM + 64 => b"000000000000000000000000", -- 0 : 
        VMEM + 65 => b"000000000000000000011001", -- 25 : 
        VMEM + 66 => b"000000000000000000000000", -- 0 : 
        VMEM + 67 => b"000000000000000000011001", -- 25 : 
        VMEM + 68 => b"000000000000000000000000", -- 0 : 
        VMEM + 69 => b"000000000000000000000000", -- 0 : 
        VMEM + 70 => b"000000000000000000000000", -- 0 : 
        VMEM + 71 => b"000000000000000000011001", -- 25 : 
        VMEM + 72 => b"000000000000000000000000", -- 0 : 
        VMEM + 73 => b"000000000000000000000000", -- 0 : 
        VMEM + 74 => b"000000000000000000000000", -- 0 : 
        VMEM + 75 => b"000000000000000000011001", -- 25 : 
        VMEM + 76 => b"000000000000000000000000", -- 0 : 
        VMEM + 77 => b"000000000000000000011001", -- 25 : 
        VMEM + 78 => b"000000000000000000000000", -- 0 : 
        VMEM + 79 => b"000000000000000000000000", -- 0 : 
        VMEM + 80 => b"000000000000000000000000", -- 0 : 
        VMEM + 81 => b"000000000000000000011001", -- 25 : 
        VMEM + 82 => b"000000000000000000011001", -- 25 : 
        VMEM + 83 => b"000000000000000000011001", -- 25 : 
        VMEM + 84 => b"000000000000000000011001", -- 25 : 
        VMEM + 85 => b"000000000000000000011001", -- 25 : 
        VMEM + 86 => b"000000000000000000000000", -- 0 : 
        VMEM + 87 => b"000000000000000000011001", -- 25 : 
        VMEM + 88 => b"000000000000000000011001", -- 25 : 
        VMEM + 89 => b"000000000000000000011001", -- 25 : 
        VMEM + 90 => b"000000000000000000000000", -- 0 : 
        VMEM + 91 => b"000000000000000000000000", -- 0 : 
        VMEM + 92 => b"000000000000000000000000", -- 0 : 
        VMEM + 93 => b"000000000000000000000000", -- 0 : 
        VMEM + 94 => b"000000000000000000000000", -- 0 : 
        VMEM + 95 => b"000000000000000000000000", -- 0 : 
        VMEM + 96 => b"000000000000000000000000", -- 0 : 
        VMEM + 97 => b"000000000000000000000000", -- 0 : 
        VMEM + 98 => b"000000000000000000000000", -- 0 : 
        VMEM + 99 => b"000000000000000000010000", -- 0 : 
        -- HEAP
        OTHERS => (OTHERS => '-')
    );

BEGIN

    -- Reading from two-port ram
    PROCESS (clk)
    BEGIN
        IF rising_edge(clk) THEN
            cpu_data_out <= p_mem(TO_INTEGER(cpu_address) + PROGRAM);
            video_data <= p_mem(TO_INTEGER(video_address) + VMEM);
        END IF;
    END PROCESS;

    -- STORE
    PROCESS (clk)
    BEGIN
        IF rising_edge(clk) THEN
            IF (cpu_we = '1') THEN
                p_mem(TO_INTEGER(cpu_address)) <= STD_LOGIC_VECTOR(cpu_data_in);
            END IF;
        END IF;
    END PROCESS;

END ARCHITECTURE;