LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY pMem IS
    PORT (
        clk : IN STD_LOGIC;
        rst: IN STD_LOGIC;
        cpu_address : IN unsigned(11 DOWNTO 0);
        cpu_data_out : OUT STD_LOGIC_VECTOR(23 DOWNTO 0);
        cpu_data_in : IN unsigned(23 DOWNTO 0);
        cpu_we : IN STD_LOGIC;
        video_address : IN unsigned(7 DOWNTO 0);
        video_data_out : OUT unsigned(6 DOWNTO 0)
    );
END pMem;

ARCHITECTURE func OF pMem IS


    TYPE p_mem_type IS ARRAY(0 TO 4095) OF STD_LOGIC_VECTOR(23 DOWNTO 0);

    CONSTANT PROGRAM : INTEGER := 0;
    CONSTANT VMEM : INTEGER := 1500;
    CONSTANT PATH : INTEGER := 1630;

    SIGNAL p_mem : p_mem_type := (
        -- PROGRAM
        PROGRAM+0 => b"01001_----_00_0_000010010001", -- start : JSR wait_for_player_input
        PROGRAM+1 => b"00000_0010_01_0_------------", -- LDI GR2, 2
        PROGRAM+2 => b"000000000000000000000010", -- 
        PROGRAM+3 => b"00001_0010_00_0_011010100101", -- ST 1700+1, GR2 // hp
        PROGRAM+4 => b"00000_0000_01_0_------------", -- LDI GR0, 34 //balloon tiletype
        PROGRAM+5 => b"000000000000000000100010", -- 
        PROGRAM+6 => b"00011_0000_01_0_------------", -- SUBI GR0, 1 //weird fix
        PROGRAM+7 => b"000000000000000000000001", -- 
        PROGRAM+8 => b"00000_0110_01_0_------------", -- push_balloon_hp : LDI GR6, 5
        PROGRAM+9 => b"000000000000000000000101", -- 
        PROGRAM+10 => b"01101_0110_--_0_------------", -- PUSH GR6
        PROGRAM+11 => b"00001_0001_11_0_010111011100", -- loop : STN 1500, GR1 // replace tiletype that was overwritten
        PROGRAM+12 => b"00001_0101_00_0_011010100100", -- ST 1700, GR5
        PROGRAM+13 => b"00000_0110_00_0_011010100100", -- LD GR6, 1700
        PROGRAM+14 => b"00011_0110_01_0_------------", -- SUBI GR6, 40
        PROGRAM+15 => b"000000000000000000101000", -- 
        PROGRAM+16 => b"01100_----_00_0_000000111101", -- BEQ player_dmg
        PROGRAM+17 => b"00001_0101_00_0_011010100100", -- new_ballon : ST 1700, GR5
        PROGRAM+18 => b"00000_0011_00_0_011010100100", -- LD GR3, 1700
        PROGRAM+19 => b"00000_0100_11_0_011001011110", -- LDN GR4, 1630 // GR4 := PATH[GR3]
        PROGRAM+20 => b"00001_0100_00_0_011010100100", -- ST 1700, GR4
        PROGRAM+21 => b"00000_0011_00_0_011010100100", -- LD GR3, 1700
        PROGRAM+22 => b"00000_0001_11_0_010111011100", -- LDN GR1, 1500 // GR1 := VMEM[GR3]
        PROGRAM+23 => b"01010_----_00_0_000001100101", -- BRA balloon_animation
        PROGRAM+24 => b"00010_0101_01_0_------------", -- check_monke : ADDI GR5, 1 // increment path index
        PROGRAM+25 => b"000000000000000000000001", -- 
        PROGRAM+26 => b"00001_0011_00_0_011010100100", -- ST 1700, GR3
        PROGRAM+27 => b"00000_0100_00_0_011010100100", -- LD GR4, 1700
        PROGRAM+28 => b"00010_0011_01_0_------------", -- ADDI GR3, 1 //right neighbour
        PROGRAM+29 => b"000000000000000000000001", -- 
        PROGRAM+30 => b"00000_0110_11_0_010111011100", -- LDN GR6, 1500
        PROGRAM+31 => b"00100_0110_01_0_------------", -- CMPI GR6, 1
        PROGRAM+32 => b"000000000000000000000001", -- 
        PROGRAM+33 => b"01100_----_00_0_000001010110", -- BEQ monke_animation
        PROGRAM+34 => b"00001_0100_00_0_011010100100", -- ST 1700, GR4
        PROGRAM+35 => b"00000_0011_00_0_011010100100", -- LD GR3, 1700
        PROGRAM+36 => b"00010_0011_01_0_------------", -- ADDI GR3, 13
        PROGRAM+37 => b"000000000000000000001101", -- 
        PROGRAM+38 => b"00000_0110_11_0_010111011100", -- LDN GR6, 1500
        PROGRAM+39 => b"00100_0110_01_0_------------", -- CMPI GR6, 1
        PROGRAM+40 => b"000000000000000000000001", -- 
        PROGRAM+41 => b"01100_----_00_0_000001010110", -- BEQ monke_animation
        PROGRAM+42 => b"00001_0100_00_0_011010100100", -- ST 1700, GR4
        PROGRAM+43 => b"00000_0011_00_0_011010100100", -- LD GR3, 1700
        PROGRAM+44 => b"00011_0011_01_0_------------", -- SUBI GR3, 1
        PROGRAM+45 => b"000000000000000000000001", -- 
        PROGRAM+46 => b"00000_0110_11_0_010111011100", -- LDN GR6, 1500
        PROGRAM+47 => b"00100_0110_01_0_------------", -- CMPI GR6, 1
        PROGRAM+48 => b"000000000000000000000001", -- 
        PROGRAM+49 => b"01100_----_00_0_000001010110", -- BEQ monke_animation
        PROGRAM+50 => b"00001_0100_00_0_011010100100", -- ST 1700, GR4
        PROGRAM+51 => b"00000_0011_00_0_011010100100", -- LD GR3, 1700
        PROGRAM+52 => b"00011_0011_01_0_------------", -- SUBI GR3, 13
        PROGRAM+53 => b"000000000000000000001101", -- 
        PROGRAM+54 => b"00000_0110_11_0_010111011100", -- LDN GR6, 1500
        PROGRAM+55 => b"00100_0110_01_0_------------", -- CMPI GR6, 1
        PROGRAM+56 => b"000000000000000000000001", -- 
        PROGRAM+57 => b"01100_----_00_0_000001010110", -- BEQ monke_animation
        PROGRAM+58 => b"00001_0100_00_0_011010100100", -- ST 1700, GR4
        PROGRAM+59 => b"00000_0011_00_0_011010100100", -- LD GR3, 1700
        PROGRAM+60 => b"01010_----_00_0_000000001011", -- BRA loop
        PROGRAM+61 => b"00000_0010_00_0_011010100101", -- player_dmg : LD GR2, 1700+1
        PROGRAM+62 => b"00011_0010_01_0_------------", -- SUBI GR2, 1
        PROGRAM+63 => b"000000000000000000000001", -- 
        PROGRAM+64 => b"00001_0010_00_0_011010100101", -- ST 1700+1, GR2
        PROGRAM+65 => b"00011_0010_01_0_------------", -- SUBI GR2, 0
        PROGRAM+66 => b"000000000000000000000000", -- 
        PROGRAM+67 => b"01100_----_00_0_000001101101", -- BEQ dead
        PROGRAM+68 => b"00000_0101_01_0_------------", -- LDI GR5, 0
        PROGRAM+69 => b"000000000000000000000000", -- 
        PROGRAM+70 => b"01010_----_00_0_000000010001", -- BRA new_ballon
        PROGRAM+71 => b"00000_0111_01_0_------------", -- balloon_dmg : LDI GR7, 1
        PROGRAM+72 => b"000000000000000000000001", -- 
        PROGRAM+73 => b"00001_0111_11_0_010111011100", -- STN 1500, GR7
        PROGRAM+74 => b"00001_0100_00_0_011010100100", -- ST 1700, GR4
        PROGRAM+75 => b"00000_0011_00_0_011010100100", -- LD GR3, 1700
        PROGRAM+76 => b"01110_0110_--_0_------------", -- POP GR6
        PROGRAM+77 => b"00011_0110_01_0_------------", -- SUBI GR6, 1  //different damage for diff monkeys?????
        PROGRAM+78 => b"000000000000000000000001", -- 
        PROGRAM+79 => b"01100_----_00_0_000001010010", -- BEQ balloon_dead
        PROGRAM+80 => b"01101_0110_--_0_------------", -- PUSH GR6
        PROGRAM+81 => b"01010_----_00_0_000000001011", -- BRA loop
        PROGRAM+82 => b"00001_0001_11_0_010111011100", -- balloon_dead : STN 1500, GR1
        PROGRAM+83 => b"00000_0101_01_0_------------", -- LDI GR5, 0
        PROGRAM+84 => b"000000000000000000000000", -- 
        PROGRAM+85 => b"01010_----_00_0_000000001000", -- BRA push_balloon_hp
        PROGRAM+86 => b"00100_0110_01_0_------------", -- monke_animation : CMPI GR6, 4
        PROGRAM+87 => b"000000000000000000000100", -- 
        PROGRAM+88 => b"01100_----_00_0_000001000111", -- BEQ balloon_dmg
        PROGRAM+89 => b"00010_0110_01_0_------------", -- ADDI GR6, 1
        PROGRAM+90 => b"000000000000000000000001", -- 
        PROGRAM+91 => b"00001_0110_11_0_010111011100", -- STN 1500, GR6
        PROGRAM+92 => b"01001_----_00_0_000010001001", -- JSR delay
        PROGRAM+93 => b"01010_----_00_0_000001010110", -- BRA monke_animation ;b
        PROGRAM+94 => b"00011_0000_01_0_------------", -- reset_anim_state : SUBI GR0, 3
        PROGRAM+95 => b"000000000000000000000011", -- 
        PROGRAM+96 => b"00001_0000_11_0_010111011100", -- STN 1500, GR0
        PROGRAM+97 => b"01001_----_00_0_000010001001", -- JSR delay
        PROGRAM+98 => b"00011_0000_01_0_------------", -- SUBI GR0, 1 ;b
        PROGRAM+99 => b"000000000000000000000001", -- 
        PROGRAM+100 => b"01010_----_00_0_000000011000", -- BRA check_monke
        PROGRAM+101 => b"00100_0000_01_0_------------", -- balloon_animation : CMPI GR0, 37
        PROGRAM+102 => b"000000000000000000100101", -- 
        PROGRAM+103 => b"01100_----_00_0_000001011110", -- BEQ reset_anim_state
        PROGRAM+104 => b"00010_0000_01_0_------------", -- ADDI GR0, 1
        PROGRAM+105 => b"000000000000000000000001", -- 
        PROGRAM+106 => b"00001_0000_11_0_010111011100", -- STN 1500, GR0
        PROGRAM+107 => b"01001_----_00_0_000010001001", -- JSR delay
        PROGRAM+108 => b"01010_----_00_0_000001100101", -- BRA balloon_animation ;b
        PROGRAM+109 => b"01010_----_00_0_000001101101", -- dead : BRA dead ;b
        PROGRAM+110 => b"00100_1111_01_1_------------", -- read_input : CMPI GR15, 1
        PROGRAM+111 => b"000000000000000000000001", -- 
        PROGRAM+112 => b"01100_----_00_0_000010010101", -- BEQ left_input // A key
        PROGRAM+113 => b"00100_1111_01_1_------------", -- CMPI GR15, 2
        PROGRAM+114 => b"000000000000000000000010", -- 
        PROGRAM+115 => b"01100_----_00_0_000010011000", -- BEQ right_input // D key
        PROGRAM+116 => b"00100_1111_01_1_------------", -- CMPI GR15, 4 // W key
        PROGRAM+117 => b"000000000000000000000100", -- 
        PROGRAM+118 => b"01100_----_00_0_000010011011", -- BEQ up_input
        PROGRAM+119 => b"00100_1111_01_1_------------", -- CMPI GR15, 8 // S key
        PROGRAM+120 => b"000000000000000000001000", -- 
        PROGRAM+121 => b"01100_----_00_0_000010011110", -- BEQ down_input
        PROGRAM+122 => b"00100_1111_01_1_------------", -- CMPI GR15, 3
        PROGRAM+123 => b"000000000000000000000011", -- 
        PROGRAM+124 => b"10000_----_--_0_------------", -- RET
        PROGRAM+125 => b"00000_1111_01_1_------------", -- mark_input_as_read : LDI GR15, 0
        PROGRAM+126 => b"000000000000000000000000", -- 
        PROGRAM+127 => b"10000_----_--_0_------------", -- RET
        PROGRAM+128 => b"00000_0000_01_0_------------", -- update_hp : LDI GR0, 54
        PROGRAM+129 => b"000000000000000000110110", -- 
        PROGRAM+130 => b"00000_0001_01_0_------------", -- LDI GR1, 11
        PROGRAM+131 => b"000000000000000000001011", -- 
        PROGRAM+132 => b"00000_0011_01_0_------------", -- LDI GR3, 4
        PROGRAM+133 => b"000000000000000000000100", -- 
        PROGRAM+134 => b"00001_0001_11_0_010111011100", -- STN 1500, GR1
        PROGRAM+135 => b"00001_0001_11_0_010111011100", -- STN 1500, GR1
        PROGRAM+136 => b"10000_----_--_0_------------", -- RET
        PROGRAM+137 => b"01101_0000_--_0_------------", -- delay : PUSH GR0
        PROGRAM+138 => b"00000_0000_01_0_------------", -- LDI GR0, 0x0FFFFF
        PROGRAM+139 => b"000011111111111111111111", -- 
        PROGRAM+140 => b"00011_0000_01_0_------------", -- delay_loop : SUBI GR0, 1
        PROGRAM+141 => b"000000000000000000000001", -- 
        PROGRAM+142 => b"01011_----_00_0_000010001100", -- BNE delay_loop
        PROGRAM+143 => b"01110_0000_--_0_------------", -- delay_end : POP GR0
        PROGRAM+144 => b"10000_----_--_0_------------", -- RET
        PROGRAM+145 => b"00100_1111_01_1_------------", -- wait_for_player_input : CMPI GR15, 3     // loop until user input
        PROGRAM+146 => b"000000000000000000000011", -- 
        PROGRAM+147 => b"01011_----_00_0_000010010001", -- BNE wait_for_player_input
        PROGRAM+148 => b"10000_----_--_0_------------", -- RET
        PROGRAM+149 => b"00000_0000_01_0_------------", -- left_input : LDI GR0, 1
        PROGRAM+150 => b"000000000000000000000001", -- 
        PROGRAM+151 => b"10000_----_--_0_------------", -- RET
        PROGRAM+152 => b"00000_0000_01_0_------------", -- right_input : LDI GR0, 2
        PROGRAM+153 => b"000000000000000000000010", -- 
        PROGRAM+154 => b"10000_----_--_0_------------", -- RET
        PROGRAM+155 => b"00000_0000_01_0_------------", -- up_input : LDI GR0, 3
        PROGRAM+156 => b"000000000000000000000011", -- 
        PROGRAM+157 => b"10000_----_--_0_------------", -- RET
        PROGRAM+158 => b"00000_0000_01_0_------------", -- down_input : LDI GR0, 4
        PROGRAM+159 => b"000000000000000000000100", -- 
        PROGRAM+160 => b"10000_----_--_0_------------", -- RET
        PROGRAM+161 => b"11111_---_--_--_------------", -- HALT
        -- VMEM
        VMEM+0 => b"000000000000000000000000", -- 0
        VMEM+1 => b"000000000000000000000000", -- 0
        VMEM+2 => b"000000000000000000000000", -- 0
        VMEM+3 => b"000000000000000000000000", -- 0
        VMEM+4 => b"000000000000000000000000", -- 0
        VMEM+5 => b"000000000000000000000000", -- 0
        VMEM+6 => b"000000000000000000000000", -- 0
        VMEM+7 => b"000000000000000000000000", -- 0
        VMEM+8 => b"000000000000000000000000", -- 0
        VMEM+9 => b"000000000000000000000000", -- 0
        VMEM+10 => b"000000000000000000110001", -- 49
        VMEM+11 => b"000000000000000000111111", -- 63
        VMEM+12 => b"000000000000000000111111", -- 63
        VMEM+13 => b"000000000000000000000000", -- 0
        VMEM+14 => b"000000000000000000011001", -- 25
        VMEM+15 => b"000000000000000000011001", -- 25
        VMEM+16 => b"000000000000000000011001", -- 25
        VMEM+17 => b"000000000000000000011001", -- 25
        VMEM+18 => b"000000000000000000011001", -- 25
        VMEM+19 => b"000000000000000000011001", -- 25
        VMEM+20 => b"000000000000000000011001", -- 25
        VMEM+21 => b"000000000000000000011001", -- 25
        VMEM+22 => b"000000000000000000000000", -- 0
        VMEM+23 => b"000000000000000000110011", -- 51
        VMEM+24 => b"000000000000000000110110", -- 54
        VMEM+25 => b"000000000000000000110110", -- 54
        VMEM+26 => b"000000000000000000000000", -- 0
        VMEM+27 => b"000000000000000000011001", -- 25
        VMEM+28 => b"000000000000000000000001", -- 1
        VMEM+29 => b"000000000000000000000000", -- 0
        VMEM+30 => b"000000000000000000000001", -- 1
        VMEM+31 => b"000000000000000000000000", -- 0
        VMEM+32 => b"000000000000000000000000", -- 0
        VMEM+33 => b"000000000000000000000000", -- 0
        VMEM+34 => b"000000000000000000011001", -- 25
        VMEM+35 => b"000000000000000000000000", -- 0
        VMEM+36 => b"000000000000000000000001", -- 1
        VMEM+37 => b"000000000000000000100110", -- 38
        VMEM+38 => b"000000000000000000000101", -- 5
        VMEM+39 => b"000000000000000000000000", -- 0
        VMEM+40 => b"000000000000000000011001", -- 25
        VMEM+41 => b"000000000000000000000000", -- 0
        VMEM+42 => b"000000000000000000011001", -- 25
        VMEM+43 => b"000000000000000000011001", -- 25
        VMEM+44 => b"000000000000000000011001", -- 25
        VMEM+45 => b"000000000000000000011001", -- 25
        VMEM+46 => b"000000000000000000011001", -- 25
        VMEM+47 => b"000000000000000000011001", -- 25
        VMEM+48 => b"000000000000000000000000", -- 0
        VMEM+49 => b"000000000000000000100110", -- 38
        VMEM+50 => b"000000000000000000100110", -- 38
        VMEM+51 => b"000000000000000000100110", -- 38
        VMEM+52 => b"000000000000000000011001", -- 25
        VMEM+53 => b"000000000000000000011001", -- 25
        VMEM+54 => b"000000000000000000000000", -- 0
        VMEM+55 => b"000000000000000000011001", -- 25
        VMEM+56 => b"000000000000000000000000", -- 0
        VMEM+57 => b"000000000000000000000000", -- 0
        VMEM+58 => b"000000000000000000000000", -- 0
        VMEM+59 => b"000000000000000000000000", -- 0
        VMEM+60 => b"000000000000000000000000", -- 0
        VMEM+61 => b"000000000000000000000000", -- 0
        VMEM+62 => b"000000000000000000001001", -- 9
        VMEM+63 => b"000000000000000000110101", -- 53
        VMEM+64 => b"000000000000000000001101", -- 13
        VMEM+65 => b"000000000000000000000000", -- 0
        VMEM+66 => b"000000000000000000000000", -- 0
        VMEM+67 => b"000000000000000000000000", -- 0
        VMEM+68 => b"000000000000000000011001", -- 25
        VMEM+69 => b"000000000000000000000000", -- 0
        VMEM+70 => b"000000000000000000011001", -- 25
        VMEM+71 => b"000000000000000000011001", -- 25
        VMEM+72 => b"000000000000000000011001", -- 25
        VMEM+73 => b"000000000000000000000000", -- 0
        VMEM+74 => b"000000000000000000000000", -- 0
        VMEM+75 => b"000000000000000000100110", -- 38
        VMEM+76 => b"000000000000000000100110", -- 38
        VMEM+77 => b"000000000000000000100110", -- 38
        VMEM+78 => b"000000000000000000000000", -- 0
        VMEM+79 => b"000000000000000000011001", -- 25
        VMEM+80 => b"000000000000000000011001", -- 25
        VMEM+81 => b"000000000000000000011001", -- 25
        VMEM+82 => b"000000000000000000000000", -- 0
        VMEM+83 => b"000000000000000000011001", -- 25
        VMEM+84 => b"000000000000000000000000", -- 0
        VMEM+85 => b"000000000000000000011001", -- 25
        VMEM+86 => b"000000000000000000000000", -- 0
        VMEM+87 => b"000000000000000000000000", -- 0
        VMEM+88 => b"000000000000000000010001", -- 17
        VMEM+89 => b"000000000000000000100110", -- 38
        VMEM+90 => b"000000000000000000010101", -- 21
        VMEM+91 => b"000000000000000000000000", -- 0
        VMEM+92 => b"000000000000000000011001", -- 25
        VMEM+93 => b"000000000000000000000000", -- 0
        VMEM+94 => b"000000000000000000000000", -- 0
        VMEM+95 => b"000000000000000000000000", -- 0
        VMEM+96 => b"000000000000000000011001", -- 25
        VMEM+97 => b"000000000000000000000000", -- 0
        VMEM+98 => b"000000000000000000011001", -- 25
        VMEM+99 => b"000000000000000000000000", -- 0
        VMEM+100 => b"000000000000000000000000", -- 0
        VMEM+101 => b"000000000000000000100110", -- 38
        VMEM+102 => b"000000000000000000100110", -- 38
        VMEM+103 => b"000000000000000000100110", -- 38
        VMEM+104 => b"000000000000000000000000", -- 0
        VMEM+105 => b"000000000000000000011001", -- 25
        VMEM+106 => b"000000000000000000011001", -- 25
        VMEM+107 => b"000000000000000000011001", -- 25
        VMEM+108 => b"000000000000000000011001", -- 25
        VMEM+109 => b"000000000000000000011001", -- 25
        VMEM+110 => b"000000000000000000000000", -- 0
        VMEM+111 => b"000000000000000000011001", -- 25
        VMEM+112 => b"000000000000000000011001", -- 25
        VMEM+113 => b"000000000000000000011001", -- 25
        VMEM+114 => b"000000000000000001000000", -- 64
        VMEM+115 => b"000000000000000001000000", -- 64
        VMEM+116 => b"000000000000000001000000", -- 64
        VMEM+117 => b"000000000000000000000000", -- 0
        VMEM+118 => b"000000000000000000000000", -- 0
        VMEM+119 => b"000000000000000000000000", -- 0
        VMEM+120 => b"000000000000000000000000", -- 0
        VMEM+121 => b"000000000000000000000000", -- 0
        VMEM+122 => b"000000000000000000000000", -- 0
        VMEM+123 => b"000000000000000000000000", -- 0
        VMEM+124 => b"000000000000000000000000", -- 0
        VMEM+125 => b"000000000000000000000000", -- 0
        VMEM+126 => b"000000000000000000000000", -- 0
        VMEM+127 => b"000000000000000000101101", -- 45
        VMEM+128 => b"000000000000000000100110", -- 38
        VMEM+129 => b"000000000000000000101111", -- 47
        -- PATH
        PATH+0 => b"000000000000000000110100", -- 52
        PATH+1 => b"000000000000000000110101", -- 53
        PATH+2 => b"000000000000000000101000", -- 40
        PATH+3 => b"000000000000000000011011", -- 27
        PATH+4 => b"000000000000000000001110", -- 14
        PATH+5 => b"000000000000000000001111", -- 15
        PATH+6 => b"000000000000000000010000", -- 16
        PATH+7 => b"000000000000000000010001", -- 17
        PATH+8 => b"000000000000000000010010", -- 18
        PATH+9 => b"000000000000000000010011", -- 19
        PATH+10 => b"000000000000000000010100", -- 20
        PATH+11 => b"000000000000000000010101", -- 21
        PATH+12 => b"000000000000000000100010", -- 34
        PATH+13 => b"000000000000000000101111", -- 47
        PATH+14 => b"000000000000000000101110", -- 46
        PATH+15 => b"000000000000000000101101", -- 45
        PATH+16 => b"000000000000000000101100", -- 44
        PATH+17 => b"000000000000000000101011", -- 43
        PATH+18 => b"000000000000000000101010", -- 42
        PATH+19 => b"000000000000000000110111", -- 55
        PATH+20 => b"000000000000000001000100", -- 68
        PATH+21 => b"000000000000000001010001", -- 81
        PATH+22 => b"000000000000000001010000", -- 80
        PATH+23 => b"000000000000000001001111", -- 79
        PATH+24 => b"000000000000000001011100", -- 92
        PATH+25 => b"000000000000000001101001", -- 105
        PATH+26 => b"000000000000000001101010", -- 106
        PATH+27 => b"000000000000000001101011", -- 107
        PATH+28 => b"000000000000000001101100", -- 108
        PATH+29 => b"000000000000000001101101", -- 109
        PATH+30 => b"000000000000000001100000", -- 96
        PATH+31 => b"000000000000000001010011", -- 83
        PATH+32 => b"000000000000000001000110", -- 70
        PATH+33 => b"000000000000000001000111", -- 71
        PATH+34 => b"000000000000000001001000", -- 72
        PATH+35 => b"000000000000000001010101", -- 85
        PATH+36 => b"000000000000000001100010", -- 98
        PATH+37 => b"000000000000000001101111", -- 111
        PATH+38 => b"000000000000000001110000", -- 112
        PATH+39 => b"000000000000000001110001", -- 113
        PATH+40 => b"000000000000000001110010", -- 114
        -- HEAP
        OTHERS => (OTHERS => '-')
    );

BEGIN

    -- Reading from two-port ram
    PROCESS (clk)
    BEGIN
        IF rising_edge(clk) THEN
            cpu_data_out <= p_mem(TO_INTEGER(cpu_address) + PROGRAM);
            video_data_out <= unsigned(p_mem(TO_INTEGER(video_address) + VMEM)(6 DOWNTO 0));
        END IF;
    END PROCESS;

    -- STORE
    PROCESS (clk)
    BEGIN
        IF rising_edge(clk) THEN
            IF (cpu_we = '1') THEN
                p_mem(TO_INTEGER(cpu_address)) <= STD_LOGIC_VECTOR(cpu_data_in);
            END IF;
        END IF;
    END PROCESS;

END ARCHITECTURE;