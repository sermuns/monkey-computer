LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY pMem IS
    PORT (
        clk : IN STD_LOGIC;
        rst: IN STD_LOGIC;
        cpu_address : IN unsigned(11 DOWNTO 0);
        cpu_data_out : OUT STD_LOGIC_VECTOR(23 DOWNTO 0);
        cpu_data_in : IN unsigned(23 DOWNTO 0);
        cpu_we : IN STD_LOGIC;
        video_address : IN unsigned(7 DOWNTO 0);
        video_data_out : OUT unsigned(6 DOWNTO 0)
    );
END pMem;

ARCHITECTURE func OF pMem IS


    TYPE p_mem_type IS ARRAY(0 TO 4095) OF STD_LOGIC_VECTOR(23 DOWNTO 0);

    CONSTANT PROGRAM : INTEGER := 0;
    CONSTANT VMEM : INTEGER := 1500;
    CONSTANT PATH : INTEGER := 1630;

    SIGNAL p_mem : p_mem_type := (
        -- PROGRAM
        PROGRAM+0 => b"00000_0000_01_0_------------", -- start : LDI GR0, 0x05FFFF
        PROGRAM+1 => b"000001011111111111111111", -- 
        PROGRAM+2 => b"00001_0000_00_0_011010101100", -- ST 1700+8, GR0
        PROGRAM+3 => b"00000_0010_01_0_------------", -- LDI GR2, 1
        PROGRAM+4 => b"000000000000000000000001", -- 
        PROGRAM+5 => b"00001_0010_00_0_011010101001", -- ST 1700+5, GR2
        PROGRAM+6 => b"00000_0010_01_0_------------", -- LDI GR2, 1
        PROGRAM+7 => b"000000000000000000000001", -- 
        PROGRAM+8 => b"00001_0010_00_0_011010100101", -- ST 1700+1, GR2 // hp
        PROGRAM+9 => b"00000_0010_01_0_------------", -- LDI GR2, 1
        PROGRAM+10 => b"000000000000000000000001", -- 
        PROGRAM+11 => b"00001_0010_00_0_011010100110", -- ST 1700+2, GR2 // hp
        PROGRAM+12 => b"00000_0010_01_0_------------", -- LDI GR2, 3
        PROGRAM+13 => b"000000000000000000000011", -- 
        PROGRAM+14 => b"00001_0010_00_0_011010100111", -- ST 1700+3, GR2 // gold
        PROGRAM+15 => b"00000_0010_01_0_------------", -- LDI GR2, 0
        PROGRAM+16 => b"000000000000000000000000", -- 
        PROGRAM+17 => b"00001_0010_00_0_011010101000", -- ST 1700+4, GR2 // gold
        PROGRAM+18 => b"01001_----_00_0_000100111000", -- JSR update_gold
        PROGRAM+19 => b"01001_----_00_0_000100101101", -- JSR update_hp
        PROGRAM+20 => b"00000_0010_01_0_------------", -- LDI GR2, 38
        PROGRAM+21 => b"000000000000000000100110", -- 
        PROGRAM+22 => b"00001_0010_00_0_011010101011", -- ST 1700+7, GR2 // save tile that cursor replaces
        PROGRAM+23 => b"00000_0010_01_0_------------", -- LDI GR2, 63
        PROGRAM+24 => b"000000000000000000111111", -- 
        PROGRAM+25 => b"00001_0010_00_0_011010101010", -- ST 1700+6, GR2 // save tile that cursor replaces
        PROGRAM+26 => b"00000_0000_01_0_------------", -- LDI GR0, 34 //balloon tiletype
        PROGRAM+27 => b"000000000000000000100010", -- 
        PROGRAM+28 => b"00011_0000_01_0_------------", -- SUBI GR0, 1 //weird fix
        PROGRAM+29 => b"000000000000000000000001", -- 
        PROGRAM+30 => b"00000_0110_00_0_011010101001", -- push_balloon_hp : LD GR6, 1700+5
        PROGRAM+31 => b"00010_0110_01_0_------------", -- ADDI GR6, 1
        PROGRAM+32 => b"000000000000000000000001", -- 
        PROGRAM+33 => b"01101_0110_--_0_------------", -- PUSH GR6
        PROGRAM+34 => b"00000_0011_00_0_011010101010", -- reset_cursor : LD GR3, 1700+6
        PROGRAM+35 => b"00000_0010_00_0_011010101011", -- LD GR2, 1700+7
        PROGRAM+36 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2 // update screen, ersätt 56 med cursorpos
        PROGRAM+37 => b"01001_----_00_0_000100001100", -- shopping_phase : JSR read_input
        PROGRAM+38 => b"00100_1000_01_0_------------", -- CMPI GR8, 1
        PROGRAM+39 => b"000000000000000000000001", -- 
        PROGRAM+40 => b"00000_1000_01_0_------------", -- LDI GR8, 0
        PROGRAM+41 => b"000000000000000000000000", -- 
        PROGRAM+42 => b"01011_----_00_0_000000100101", -- BNE shopping_phase // continue shopping
        PROGRAM+43 => b"01010_----_00_0_000000101101", -- BRA loop
        PROGRAM+44 => b"00001_0001_11_0_010111011100", -- pre_loop : STN 1500, GR1 // replace tiletype that was overwritten
        PROGRAM+45 => b"01101_0101_--_0_------------", -- loop : PUSH GR5
        PROGRAM+46 => b"01110_0110_--_0_------------", -- POP GR6
        PROGRAM+47 => b"00011_0110_01_0_------------", -- SUBI GR6, 40 // 40 is the end of the map! taken from path index.
        PROGRAM+48 => b"000000000000000000101000", -- 
        PROGRAM+49 => b"01100_----_00_0_000010011010", -- BEQ player_dmg
        PROGRAM+50 => b"01101_0101_--_0_------------", -- new_ballon : PUSH GR5
        PROGRAM+51 => b"01110_0011_--_0_------------", -- POP GR3
        PROGRAM+52 => b"00000_0100_11_0_011001011110", -- LDN GR4, 1630 // GR4 := PATH[GR3]
        PROGRAM+53 => b"01101_0100_--_0_------------", -- PUSH GR4
        PROGRAM+54 => b"01110_0011_--_0_------------", -- POP GR3
        PROGRAM+55 => b"00000_0001_11_0_010111011100", -- LDN GR1, 1500 // GR1 := VMEM[GR3]
        PROGRAM+56 => b"01010_----_00_0_000011100011", -- BRA balloon_animation
        PROGRAM+57 => b"00010_0101_01_0_------------", -- check_monke : ADDI GR5, 1 // increment path index
        PROGRAM+58 => b"000000000000000000000001", -- 
        PROGRAM+59 => b"01101_0011_--_0_------------", -- PUSH GR3
        PROGRAM+60 => b"01110_0100_--_0_------------", -- POP GR4
        PROGRAM+61 => b"00010_0011_01_0_------------", -- ADDI GR3, 1 //right neighbour
        PROGRAM+62 => b"000000000000000000000001", -- 
        PROGRAM+63 => b"00000_0110_11_0_010111011100", -- LDN GR6, 1500
        PROGRAM+64 => b"00100_0110_01_0_------------", -- CMPI GR6, 1
        PROGRAM+65 => b"000000000000000000000001", -- 
        PROGRAM+66 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+67 => b"00100_0110_01_0_------------", -- CMPI GR6, 5
        PROGRAM+68 => b"000000000000000000000101", -- 
        PROGRAM+69 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+70 => b"00100_0110_01_0_------------", -- CMPI GR6, 9
        PROGRAM+71 => b"000000000000000000001001", -- 
        PROGRAM+72 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+73 => b"00100_0110_01_0_------------", -- CMPI GR6, 13
        PROGRAM+74 => b"000000000000000000001101", -- 
        PROGRAM+75 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+76 => b"00100_0110_01_0_------------", -- CMPI GR6, 17
        PROGRAM+77 => b"000000000000000000010001", -- 
        PROGRAM+78 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+79 => b"00100_0110_01_0_------------", -- CMPI GR6, 21
        PROGRAM+80 => b"000000000000000000010101", -- 
        PROGRAM+81 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+82 => b"01101_0100_--_0_------------", -- PUSH GR4
        PROGRAM+83 => b"01110_0011_--_0_------------", -- POP GR3
        PROGRAM+84 => b"00010_0011_01_0_------------", -- ADDI GR3, 13
        PROGRAM+85 => b"000000000000000000001101", -- 
        PROGRAM+86 => b"00000_0110_11_0_010111011100", -- LDN GR6, 1500
        PROGRAM+87 => b"00100_0110_01_0_------------", -- CMPI GR6, 1
        PROGRAM+88 => b"000000000000000000000001", -- 
        PROGRAM+89 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+90 => b"00100_0110_01_0_------------", -- CMPI GR6, 5
        PROGRAM+91 => b"000000000000000000000101", -- 
        PROGRAM+92 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+93 => b"00100_0110_01_0_------------", -- CMPI GR6, 9
        PROGRAM+94 => b"000000000000000000001001", -- 
        PROGRAM+95 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+96 => b"00100_0110_01_0_------------", -- CMPI GR6, 13
        PROGRAM+97 => b"000000000000000000001101", -- 
        PROGRAM+98 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+99 => b"00100_0110_01_0_------------", -- CMPI GR6, 17
        PROGRAM+100 => b"000000000000000000010001", -- 
        PROGRAM+101 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+102 => b"00100_0110_01_0_------------", -- CMPI GR6, 21
        PROGRAM+103 => b"000000000000000000010101", -- 
        PROGRAM+104 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+105 => b"01101_0100_--_0_------------", -- PUSH GR4
        PROGRAM+106 => b"01110_0011_--_0_------------", -- POP GR3
        PROGRAM+107 => b"00011_0011_01_0_------------", -- SUBI GR3, 1
        PROGRAM+108 => b"000000000000000000000001", -- 
        PROGRAM+109 => b"00000_0110_11_0_010111011100", -- LDN GR6, 1500
        PROGRAM+110 => b"00100_0110_01_0_------------", -- CMPI GR6, 1
        PROGRAM+111 => b"000000000000000000000001", -- 
        PROGRAM+112 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+113 => b"00100_0110_01_0_------------", -- CMPI GR6, 5
        PROGRAM+114 => b"000000000000000000000101", -- 
        PROGRAM+115 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+116 => b"00100_0110_01_0_------------", -- CMPI GR6, 9
        PROGRAM+117 => b"000000000000000000001001", -- 
        PROGRAM+118 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+119 => b"00100_0110_01_0_------------", -- CMPI GR6, 13
        PROGRAM+120 => b"000000000000000000001101", -- 
        PROGRAM+121 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+122 => b"00100_0110_01_0_------------", -- CMPI GR6, 17
        PROGRAM+123 => b"000000000000000000010001", -- 
        PROGRAM+124 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+125 => b"00100_0110_01_0_------------", -- CMPI GR6, 21
        PROGRAM+126 => b"000000000000000000010101", -- 
        PROGRAM+127 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+128 => b"01101_0100_--_0_------------", -- PUSH GR4
        PROGRAM+129 => b"01110_0011_--_0_------------", -- POP GR3
        PROGRAM+130 => b"00011_0011_01_0_------------", -- SUBI GR3, 13
        PROGRAM+131 => b"000000000000000000001101", -- 
        PROGRAM+132 => b"00000_0110_11_0_010111011100", -- LDN GR6, 1500
        PROGRAM+133 => b"00100_0110_01_0_------------", -- CMPI GR6, 1
        PROGRAM+134 => b"000000000000000000000001", -- 
        PROGRAM+135 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+136 => b"00100_0110_01_0_------------", -- CMPI GR6, 5
        PROGRAM+137 => b"000000000000000000000101", -- 
        PROGRAM+138 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+139 => b"00100_0110_01_0_------------", -- CMPI GR6, 9
        PROGRAM+140 => b"000000000000000000001001", -- 
        PROGRAM+141 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+142 => b"00100_0110_01_0_------------", -- CMPI GR6, 13
        PROGRAM+143 => b"000000000000000000001101", -- 
        PROGRAM+144 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+145 => b"00100_0110_01_0_------------", -- CMPI GR6, 17
        PROGRAM+146 => b"000000000000000000010001", -- 
        PROGRAM+147 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+148 => b"00100_0110_01_0_------------", -- CMPI GR6, 21
        PROGRAM+149 => b"000000000000000000010101", -- 
        PROGRAM+150 => b"01100_----_00_0_000011000101", -- BEQ monke_animation
        PROGRAM+151 => b"01101_0100_--_0_------------", -- PUSH GR4
        PROGRAM+152 => b"01110_0011_--_0_------------", -- POP GR3
        PROGRAM+153 => b"01010_----_00_0_000000101100", -- BRA pre_loop
        PROGRAM+154 => b"00000_0010_00_0_011010100101", -- player_dmg : LD GR2, 1700+1
        PROGRAM+155 => b"00100_0010_01_0_------------", -- CMPI GR2, 0
        PROGRAM+156 => b"000000000000000000000000", -- 
        PROGRAM+157 => b"01100_----_00_0_001011001000", -- BEQ decrement_of_hp
        PROGRAM+158 => b"00011_0010_01_0_------------", -- SUBI GR2, 1
        PROGRAM+159 => b"000000000000000000000001", -- 
        PROGRAM+160 => b"00001_0010_00_0_011010100101", -- ST 1700+1, GR2
        PROGRAM+161 => b"01001_----_00_0_000100101101", -- player_dmg_2 : JSR update_hp
        PROGRAM+162 => b"00000_0010_00_0_011010100101", -- LD GR2, 1700+1
        PROGRAM+163 => b"00010_0010_00_0_011010100110", -- ADD GR2, 1700+2
        PROGRAM+164 => b"01100_----_00_0_000011110001", -- BEQ dead
        PROGRAM+165 => b"00000_0101_01_0_------------", -- LDI GR5, 0
        PROGRAM+166 => b"000000000000000000000000", -- 
        PROGRAM+167 => b"01010_----_00_0_000000110010", -- BRA new_ballon
        PROGRAM+168 => b"00011_0110_01_0_------------", -- balloon_dmg : SUBI GR6, 3
        PROGRAM+169 => b"000000000000000000000011", -- 
        PROGRAM+170 => b"00001_0110_11_0_010111011100", -- STN 1500, GR6
        PROGRAM+171 => b"01101_0100_--_0_------------", -- PUSH GR4
        PROGRAM+172 => b"01110_0011_--_0_------------", -- POP GR3
        PROGRAM+173 => b"01110_0110_--_0_------------", -- POP GR6
        PROGRAM+174 => b"00011_0110_01_0_------------", -- SUBI GR6, 1  //different damage for diff monkeys?????
        PROGRAM+175 => b"000000000000000000000001", -- 
        PROGRAM+176 => b"01100_----_00_0_000010110011", -- BEQ balloon_dead
        PROGRAM+177 => b"01101_0110_--_0_------------", -- PUSH GR6
        PROGRAM+178 => b"01010_----_00_0_000000101100", -- BRA pre_loop
        PROGRAM+179 => b"01101_0011_--_0_------------", -- balloon_dead : PUSH GR3
        PROGRAM+180 => b"00001_0001_11_0_010111011100", -- STN 1500, GR1
        PROGRAM+181 => b"00000_0101_01_0_------------", -- LDI GR5, 0
        PROGRAM+182 => b"000000000000000000000000", -- 
        PROGRAM+183 => b"00000_0111_00_0_011010100111", -- LD GR7, 1700+3
        PROGRAM+184 => b"00010_0111_01_0_------------", -- ADDI GR7, 1 // current gold reward.
        PROGRAM+185 => b"000000000000000000000001", -- 
        PROGRAM+186 => b"00100_0111_01_0_------------", -- CMPI GR7, 10
        PROGRAM+187 => b"000000000000000000001010", -- 
        PROGRAM+188 => b"01100_----_00_0_001010110100", -- BEQ increment_of_gold
        PROGRAM+189 => b"00001_0111_00_0_011010100111", -- ST 1700+3, GR7
        PROGRAM+190 => b"01001_----_00_0_000100111000", -- balloon_dead2 : JSR update_gold
        PROGRAM+191 => b"00000_0011_00_0_011010101001", -- LD GR3, 1700+5
        PROGRAM+192 => b"00010_0011_01_0_------------", -- ADDI GR3, 1
        PROGRAM+193 => b"000000000000000000000001", -- 
        PROGRAM+194 => b"00001_0011_00_0_011010101001", -- ST 1700+5, GR3
        PROGRAM+195 => b"01110_0011_--_0_------------", -- POP GR3
        PROGRAM+196 => b"01010_----_00_0_000000011110", -- BRA push_balloon_hp
        PROGRAM+197 => b"00100_0110_01_0_------------", -- monke_animation : CMPI GR6, 4
        PROGRAM+198 => b"000000000000000000000100", -- 
        PROGRAM+199 => b"01100_----_00_0_000010101000", -- BEQ balloon_dmg
        PROGRAM+200 => b"00100_0110_01_0_------------", -- CMPI GR6, 8
        PROGRAM+201 => b"000000000000000000001000", -- 
        PROGRAM+202 => b"01100_----_00_0_000010101000", -- BEQ balloon_dmg
        PROGRAM+203 => b"00100_0110_01_0_------------", -- CMPI GR6, 12
        PROGRAM+204 => b"000000000000000000001100", -- 
        PROGRAM+205 => b"01100_----_00_0_000010101000", -- BEQ balloon_dmg
        PROGRAM+206 => b"00100_0110_01_0_------------", -- CMPI GR6, 16
        PROGRAM+207 => b"000000000000000000010000", -- 
        PROGRAM+208 => b"01100_----_00_0_000010101000", -- BEQ balloon_dmg
        PROGRAM+209 => b"00100_0110_01_0_------------", -- CMPI GR6, 20
        PROGRAM+210 => b"000000000000000000010100", -- 
        PROGRAM+211 => b"01100_----_00_0_000010101000", -- BEQ balloon_dmg
        PROGRAM+212 => b"00100_0110_01_0_------------", -- CMPI GR6, 24
        PROGRAM+213 => b"000000000000000000011000", -- 
        PROGRAM+214 => b"01100_----_00_0_000010101000", -- BEQ balloon_dmg
        PROGRAM+215 => b"00010_0110_01_0_------------", -- ADDI GR6, 1
        PROGRAM+216 => b"000000000000000000000001", -- 
        PROGRAM+217 => b"00001_0110_11_0_010111011100", -- STN 1500, GR6
        PROGRAM+218 => b"01001_----_00_0_001011010100", -- JSR delay
        PROGRAM+219 => b"01010_----_00_0_000011000101", -- BRA monke_animation ;b
        PROGRAM+220 => b"00011_0000_01_0_------------", -- reset_anim_state : SUBI GR0, 3
        PROGRAM+221 => b"000000000000000000000011", -- 
        PROGRAM+222 => b"00001_0000_11_0_010111011100", -- STN 1500, GR0
        PROGRAM+223 => b"01001_----_00_0_001011010100", -- JSR delay
        PROGRAM+224 => b"00011_0000_01_0_------------", -- SUBI GR0, 1 ;b
        PROGRAM+225 => b"000000000000000000000001", -- 
        PROGRAM+226 => b"01010_----_00_0_000000111001", -- BRA check_monke
        PROGRAM+227 => b"00010_0000_01_0_------------", -- balloon_animation : ADDI GR0, 1
        PROGRAM+228 => b"000000000000000000000001", -- 
        PROGRAM+229 => b"00100_0000_01_0_------------", -- CMPI GR0, 29
        PROGRAM+230 => b"000000000000000000011101", -- 
        PROGRAM+231 => b"01100_----_00_0_000011011100", -- BEQ reset_anim_state
        PROGRAM+232 => b"00100_0000_01_0_------------", -- CMPI GR0, 33
        PROGRAM+233 => b"000000000000000000100001", -- 
        PROGRAM+234 => b"01100_----_00_0_000011011100", -- BEQ reset_anim_state
        PROGRAM+235 => b"00100_0000_01_0_------------", -- CMPI GR0, 37
        PROGRAM+236 => b"000000000000000000100101", -- 
        PROGRAM+237 => b"01100_----_00_0_000011011100", -- BEQ reset_anim_state
        PROGRAM+238 => b"00001_0000_11_0_010111011100", -- STN 1500, GR0
        PROGRAM+239 => b"01001_----_00_0_001011010100", -- JSR delay
        PROGRAM+240 => b"01010_----_00_0_000011100011", -- BRA balloon_animation ;b
        PROGRAM+241 => b"11111_----_--_0_------------", -- dead : HALT
        PROGRAM+242 => b"00100_1111_01_1_------------", -- wait_for_break : CMPI GR15, 0b11111
        PROGRAM+243 => b"000000000000000000011111", -- 
        PROGRAM+244 => b"01011_----_00_0_000011110010", -- BNE wait_for_break
        PROGRAM+245 => b"10000_----_--_0_------------", -- RET
        PROGRAM+246 => b"00100_1111_01_1_------------", -- wait_until_break_is_gone : CMPI GR15, 0b11111
        PROGRAM+247 => b"000000000000000000011111", -- 
        PROGRAM+248 => b"01100_----_00_0_000011110110", -- BEQ wait_until_break_is_gone
        PROGRAM+249 => b"10000_----_--_0_------------", -- RET
        PROGRAM+250 => b"01101_0000_--_0_------------", -- low_delay : PUSH GR0
        PROGRAM+251 => b"00000_0000_01_0_------------", -- LDI GR0, 0x00FFFF
        PROGRAM+252 => b"000000001111111111111111", -- 
        PROGRAM+253 => b"00001_0000_00_0_011010101100", -- ST 1700+8, GR0
        PROGRAM+254 => b"01110_0000_--_0_------------", -- POP GR0
        PROGRAM+255 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+256 => b"01101_0000_--_0_------------", -- mid_delay : PUSH GR0
        PROGRAM+257 => b"00000_0000_01_0_------------", -- LDI GR0, 0x05FFFF
        PROGRAM+258 => b"000001011111111111111111", -- 
        PROGRAM+259 => b"00001_0000_00_0_011010101100", -- ST 1700+8, GR0
        PROGRAM+260 => b"01110_0000_--_0_------------", -- POP GR0
        PROGRAM+261 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+262 => b"01101_0000_--_0_------------", -- high_delay : PUSH GR0
        PROGRAM+263 => b"00000_0000_01_0_------------", -- LDI GR0, 0x0FFFFF
        PROGRAM+264 => b"000011111111111111111111", -- 
        PROGRAM+265 => b"00001_0000_00_0_011010101100", -- ST 1700+8, GR0
        PROGRAM+266 => b"01110_0000_--_0_------------", -- POP GR0
        PROGRAM+267 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+268 => b"01001_----_00_0_000011110010", -- read_input : JSR wait_for_break
        PROGRAM+269 => b"01001_----_00_0_000011110110", -- JSR wait_until_break_is_gone
        PROGRAM+270 => b"00100_1111_01_1_------------", -- CMPI GR15, 0b10001
        PROGRAM+271 => b"000000000000000000010001", -- 
        PROGRAM+272 => b"01100_----_00_0_000011111010", -- BEQ low_delay
        PROGRAM+273 => b"00100_1111_01_1_------------", -- CMPI GR15, 0b10010
        PROGRAM+274 => b"000000000000000000010010", -- 
        PROGRAM+275 => b"01100_----_00_0_000100000000", -- BEQ mid_delay
        PROGRAM+276 => b"00100_1111_01_1_------------", -- CMPI GR15, 0b10011
        PROGRAM+277 => b"000000000000000000010011", -- 
        PROGRAM+278 => b"01100_----_00_0_000100000110", -- BEQ high_delay
        PROGRAM+279 => b"00100_1111_01_1_------------", -- CMPI GR15, 1
        PROGRAM+280 => b"000000000000000000000001", -- 
        PROGRAM+281 => b"01100_----_00_0_000101000011", -- BEQ left_input // A key
        PROGRAM+282 => b"00100_1111_01_1_------------", -- CMPI GR15, 2
        PROGRAM+283 => b"000000000000000000000010", -- 
        PROGRAM+284 => b"01100_----_00_0_000101110101", -- BEQ right_input // D key
        PROGRAM+285 => b"00100_1111_01_1_------------", -- CMPI GR15, 4 // W key
        PROGRAM+286 => b"000000000000000000000100", -- 
        PROGRAM+287 => b"01100_----_00_0_000110100111", -- BEQ up_input
        PROGRAM+288 => b"00100_1111_01_1_------------", -- CMPI GR15, 8 // S key
        PROGRAM+289 => b"000000000000000000001000", -- 
        PROGRAM+290 => b"01100_----_00_0_000111011001", -- BEQ down_input
        PROGRAM+291 => b"00100_1111_01_1_------------", -- CMPI GR15, 3 // Space
        PROGRAM+292 => b"000000000000000000000011", -- 
        PROGRAM+293 => b"01100_----_00_0_001000001011", -- BEQ confirm_input_pick
        PROGRAM+294 => b"00100_1111_01_1_------------", -- CMPI GR15, 5 // Enter key
        PROGRAM+295 => b"000000000000000000000101", -- 
        PROGRAM+296 => b"01100_----_00_0_001010101110", -- BEQ continue_game
        PROGRAM+297 => b"10000_----_--_0_------------", -- RET
        PROGRAM+298 => b"00000_1111_01_1_------------", -- read_input_end : LDI GR15, 0
        PROGRAM+299 => b"000000000000000000000000", -- 
        PROGRAM+300 => b"10000_----_--_0_------------", -- RET
        PROGRAM+301 => b"01101_0010_--_0_------------", -- update_hp : PUSH GR2
        PROGRAM+302 => b"00000_0010_00_0_011010100101", -- LD GR2, 1700+1
        PROGRAM+303 => b"00010_0010_01_0_------------", -- ADDI GR2, 54
        PROGRAM+304 => b"000000000000000000110110", -- 
        PROGRAM+305 => b"00001_0010_00_0_010111101000", -- ST 1500+12, GR2
        PROGRAM+306 => b"00000_0010_00_0_011010100110", -- LD GR2, 1700+2
        PROGRAM+307 => b"00010_0010_01_0_------------", -- ADDI GR2, 54
        PROGRAM+308 => b"000000000000000000110110", -- 
        PROGRAM+309 => b"00001_0010_00_0_010111100111", -- ST 1500+11, GR2
        PROGRAM+310 => b"01110_0010_--_0_------------", -- POP GR2
        PROGRAM+311 => b"10000_----_--_0_------------", -- RET
        PROGRAM+312 => b"01101_0010_--_0_------------", -- update_gold : PUSH GR2
        PROGRAM+313 => b"00000_0010_00_0_011010100111", -- LD GR2, 1700+3
        PROGRAM+314 => b"00010_0010_01_0_------------", -- ADDI GR2, 54
        PROGRAM+315 => b"000000000000000000110110", -- 
        PROGRAM+316 => b"00001_0010_00_0_010111110101", -- ST 1500+25, GR2
        PROGRAM+317 => b"00000_0010_00_0_011010101000", -- LD GR2, 1700+4
        PROGRAM+318 => b"00010_0010_01_0_------------", -- ADDI GR2, 54
        PROGRAM+319 => b"000000000000000000110110", -- 
        PROGRAM+320 => b"00001_0010_00_0_010111110100", -- ST 1500+24, GR2
        PROGRAM+321 => b"01110_0010_--_0_------------", -- POP GR2
        PROGRAM+322 => b"10000_----_--_0_------------", -- RET
        PROGRAM+323 => b"00000_0010_00_0_011010101011", -- left_input : LD GR2, 1700+7
        PROGRAM+324 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+325 => b"00001_0010_11_0_010111011100", -- STN 1500,GR2
        PROGRAM+326 => b"00011_0011_01_0_------------", -- SUBI GR3, 1
        PROGRAM+327 => b"000000000000000000000001", -- 
        PROGRAM+328 => b"00001_0011_00_0_011010101010", -- ST 1700+6, GR3
        PROGRAM+329 => b"00000_0010_11_0_010111011100", -- LDN GR2, 1500
        PROGRAM+330 => b"00001_0010_00_0_011010101011", -- ST 1700+7, GR2
        PROGRAM+331 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+332 => b"00000_0010_00_0_011010101011", -- LD GR2, 1700+7
        PROGRAM+333 => b"00100_0010_01_0_------------", -- CMPI GR2, 0
        PROGRAM+334 => b"000000000000000000000000", -- 
        PROGRAM+335 => b"01100_----_00_0_001011100001", -- BEQ set_highlighted_grass
        PROGRAM+336 => b"00100_0010_01_0_------------", -- CMPI GR2, 1
        PROGRAM+337 => b"000000000000000000000001", -- 
        PROGRAM+338 => b"01100_----_00_0_001011111001", -- BEQ set_highlighted_monkey1
        PROGRAM+339 => b"00100_0010_01_0_------------", -- CMPI GR2, 5
        PROGRAM+340 => b"000000000000000000000101", -- 
        PROGRAM+341 => b"01100_----_00_0_001011111101", -- BEQ set_highlighted_monkey2
        PROGRAM+342 => b"00100_0010_01_0_------------", -- CMPI GR2, 9
        PROGRAM+343 => b"000000000000000000001001", -- 
        PROGRAM+344 => b"01100_----_00_0_001100000001", -- BEQ set_highlighted_monkey3
        PROGRAM+345 => b"00100_0010_01_0_------------", -- CMPI GR2, 13
        PROGRAM+346 => b"000000000000000000001101", -- 
        PROGRAM+347 => b"01100_----_00_0_001100000101", -- BEQ set_highlighted_monkey4
        PROGRAM+348 => b"00100_0010_01_0_------------", -- CMPI GR2, 17
        PROGRAM+349 => b"000000000000000000010001", -- 
        PROGRAM+350 => b"01100_----_00_0_001100001001", -- BEQ set_highlighted_monkey5
        PROGRAM+351 => b"00100_0010_01_0_------------", -- CMPI GR2, 21
        PROGRAM+352 => b"000000000000000000010101", -- 
        PROGRAM+353 => b"01100_----_00_0_001100001101", -- BEQ set_highlighted_monkey6
        PROGRAM+354 => b"00100_0010_01_0_------------", -- CMPI GR2, 25
        PROGRAM+355 => b"000000000000000000011001", -- 
        PROGRAM+356 => b"01100_----_00_0_001011100101", -- BEQ set_highlighted_path
        PROGRAM+357 => b"00100_0010_01_0_------------", -- CMPI GR2, 38
        PROGRAM+358 => b"000000000000000000100110", -- 
        PROGRAM+359 => b"01100_----_00_0_001011101101", -- BEQ set_highlighted_black
        PROGRAM+360 => b"00100_0010_01_0_------------", -- CMPI GR2, 45
        PROGRAM+361 => b"000000000000000000101101", -- 
        PROGRAM+362 => b"01100_----_00_0_001011110001", -- BEQ set_highlighted_reset
        PROGRAM+363 => b"00100_0010_01_0_------------", -- CMPI GR2, 47
        PROGRAM+364 => b"000000000000000000101111", -- 
        PROGRAM+365 => b"01100_----_00_0_001011110101", -- BEQ set_highlighted_quit
        PROGRAM+366 => b"00100_0010_01_0_------------", -- CMPI GR2, 50
        PROGRAM+367 => b"000000000000000000110010", -- 
        PROGRAM+368 => b"01100_----_00_0_001011101001", -- BEQ set_highlighted_continue
        PROGRAM+369 => b"00000_0010_01_0_------------", -- LDI GR2, 53
        PROGRAM+370 => b"000000000000000000110101", -- 
        PROGRAM+371 => b"00001_0010_11_0_010111011100", -- STN 1500,GR2
        PROGRAM+372 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+373 => b"00000_0010_00_0_011010101011", -- right_input : LD GR2, 1700+7
        PROGRAM+374 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+375 => b"00001_0010_11_0_010111011100", -- STN 1500,GR2
        PROGRAM+376 => b"00010_0011_01_0_------------", -- ADDI GR3, 1
        PROGRAM+377 => b"000000000000000000000001", -- 
        PROGRAM+378 => b"00001_0011_00_0_011010101010", -- ST 1700+6, GR3
        PROGRAM+379 => b"00000_0010_11_0_010111011100", -- LDN GR2, 1500
        PROGRAM+380 => b"00001_0010_00_0_011010101011", -- ST 1700+7, GR2
        PROGRAM+381 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+382 => b"00000_0010_00_0_011010101011", -- LD GR2, 1700+7
        PROGRAM+383 => b"00100_0010_01_0_------------", -- CMPI GR2, 0
        PROGRAM+384 => b"000000000000000000000000", -- 
        PROGRAM+385 => b"01100_----_00_0_001011100001", -- BEQ set_highlighted_grass
        PROGRAM+386 => b"00100_0010_01_0_------------", -- CMPI GR2, 1
        PROGRAM+387 => b"000000000000000000000001", -- 
        PROGRAM+388 => b"01100_----_00_0_001011111001", -- BEQ set_highlighted_monkey1
        PROGRAM+389 => b"00100_0010_01_0_------------", -- CMPI GR2, 5
        PROGRAM+390 => b"000000000000000000000101", -- 
        PROGRAM+391 => b"01100_----_00_0_001011111101", -- BEQ set_highlighted_monkey2
        PROGRAM+392 => b"00100_0010_01_0_------------", -- CMPI GR2, 9
        PROGRAM+393 => b"000000000000000000001001", -- 
        PROGRAM+394 => b"01100_----_00_0_001100000001", -- BEQ set_highlighted_monkey3
        PROGRAM+395 => b"00100_0010_01_0_------------", -- CMPI GR2, 13
        PROGRAM+396 => b"000000000000000000001101", -- 
        PROGRAM+397 => b"01100_----_00_0_001100000101", -- BEQ set_highlighted_monkey4
        PROGRAM+398 => b"00100_0010_01_0_------------", -- CMPI GR2, 17
        PROGRAM+399 => b"000000000000000000010001", -- 
        PROGRAM+400 => b"01100_----_00_0_001100001001", -- BEQ set_highlighted_monkey5
        PROGRAM+401 => b"00100_0010_01_0_------------", -- CMPI GR2, 21
        PROGRAM+402 => b"000000000000000000010101", -- 
        PROGRAM+403 => b"01100_----_00_0_001100001101", -- BEQ set_highlighted_monkey6
        PROGRAM+404 => b"00100_0010_01_0_------------", -- CMPI GR2, 25
        PROGRAM+405 => b"000000000000000000011001", -- 
        PROGRAM+406 => b"01100_----_00_0_001011100101", -- BEQ set_highlighted_path
        PROGRAM+407 => b"00100_0010_01_0_------------", -- CMPI GR2, 38
        PROGRAM+408 => b"000000000000000000100110", -- 
        PROGRAM+409 => b"01100_----_00_0_001011101101", -- BEQ set_highlighted_black
        PROGRAM+410 => b"00100_0010_01_0_------------", -- CMPI GR2, 45
        PROGRAM+411 => b"000000000000000000101101", -- 
        PROGRAM+412 => b"01100_----_00_0_001011110001", -- BEQ set_highlighted_reset
        PROGRAM+413 => b"00100_0010_01_0_------------", -- CMPI GR2, 47
        PROGRAM+414 => b"000000000000000000101111", -- 
        PROGRAM+415 => b"01100_----_00_0_001011110101", -- BEQ set_highlighted_quit
        PROGRAM+416 => b"00100_0010_01_0_------------", -- CMPI GR2, 50
        PROGRAM+417 => b"000000000000000000110010", -- 
        PROGRAM+418 => b"01100_----_00_0_001011101001", -- BEQ set_highlighted_continue
        PROGRAM+419 => b"00000_0010_01_0_------------", -- LDI GR2, 53
        PROGRAM+420 => b"000000000000000000110101", -- 
        PROGRAM+421 => b"00001_0010_11_0_010111011100", -- STN 1500,GR2
        PROGRAM+422 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+423 => b"00000_0010_00_0_011010101011", -- up_input : LD GR2, 1700+7
        PROGRAM+424 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+425 => b"00001_0010_11_0_010111011100", -- STN 1500,GR2
        PROGRAM+426 => b"00011_0011_01_0_------------", -- SUBI GR3, 13
        PROGRAM+427 => b"000000000000000000001101", -- 
        PROGRAM+428 => b"00001_0011_00_0_011010101010", -- ST 1700+6, GR3
        PROGRAM+429 => b"00000_0010_11_0_010111011100", -- LDN GR2, 1500
        PROGRAM+430 => b"00001_0010_00_0_011010101011", -- ST 1700+7, GR2
        PROGRAM+431 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+432 => b"00000_0010_00_0_011010101011", -- LD GR2, 1700+7
        PROGRAM+433 => b"00100_0010_01_0_------------", -- CMPI GR2, 0
        PROGRAM+434 => b"000000000000000000000000", -- 
        PROGRAM+435 => b"01100_----_00_0_001011100001", -- BEQ set_highlighted_grass
        PROGRAM+436 => b"00100_0010_01_0_------------", -- CMPI GR2, 1
        PROGRAM+437 => b"000000000000000000000001", -- 
        PROGRAM+438 => b"01100_----_00_0_001011111001", -- BEQ set_highlighted_monkey1
        PROGRAM+439 => b"00100_0010_01_0_------------", -- CMPI GR2, 5
        PROGRAM+440 => b"000000000000000000000101", -- 
        PROGRAM+441 => b"01100_----_00_0_001011111101", -- BEQ set_highlighted_monkey2
        PROGRAM+442 => b"00100_0010_01_0_------------", -- CMPI GR2, 9
        PROGRAM+443 => b"000000000000000000001001", -- 
        PROGRAM+444 => b"01100_----_00_0_001100000001", -- BEQ set_highlighted_monkey3
        PROGRAM+445 => b"00100_0010_01_0_------------", -- CMPI GR2, 13
        PROGRAM+446 => b"000000000000000000001101", -- 
        PROGRAM+447 => b"01100_----_00_0_001100000101", -- BEQ set_highlighted_monkey4
        PROGRAM+448 => b"00100_0010_01_0_------------", -- CMPI GR2, 17
        PROGRAM+449 => b"000000000000000000010001", -- 
        PROGRAM+450 => b"01100_----_00_0_001100001001", -- BEQ set_highlighted_monkey5
        PROGRAM+451 => b"00100_0010_01_0_------------", -- CMPI GR2, 21
        PROGRAM+452 => b"000000000000000000010101", -- 
        PROGRAM+453 => b"01100_----_00_0_001100001101", -- BEQ set_highlighted_monkey6
        PROGRAM+454 => b"00100_0010_01_0_------------", -- CMPI GR2, 25
        PROGRAM+455 => b"000000000000000000011001", -- 
        PROGRAM+456 => b"01100_----_00_0_001011100101", -- BEQ set_highlighted_path
        PROGRAM+457 => b"00100_0010_01_0_------------", -- CMPI GR2, 38
        PROGRAM+458 => b"000000000000000000100110", -- 
        PROGRAM+459 => b"01100_----_00_0_001011101101", -- BEQ set_highlighted_black
        PROGRAM+460 => b"00100_0010_01_0_------------", -- CMPI GR2, 45
        PROGRAM+461 => b"000000000000000000101101", -- 
        PROGRAM+462 => b"01100_----_00_0_001011110001", -- BEQ set_highlighted_reset
        PROGRAM+463 => b"00100_0010_01_0_------------", -- CMPI GR2, 47
        PROGRAM+464 => b"000000000000000000101111", -- 
        PROGRAM+465 => b"01100_----_00_0_001011110101", -- BEQ set_highlighted_quit
        PROGRAM+466 => b"00100_0010_01_0_------------", -- CMPI GR2, 50
        PROGRAM+467 => b"000000000000000000110010", -- 
        PROGRAM+468 => b"01100_----_00_0_001011101001", -- BEQ set_highlighted_continue
        PROGRAM+469 => b"00000_0010_01_0_------------", -- LDI GR2, 53
        PROGRAM+470 => b"000000000000000000110101", -- 
        PROGRAM+471 => b"00001_0010_11_0_010111011100", -- STN 1500,GR2
        PROGRAM+472 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+473 => b"00000_0010_00_0_011010101011", -- down_input : LD GR2, 1700+7
        PROGRAM+474 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+475 => b"00001_0010_11_0_010111011100", -- STN 1500,GR2
        PROGRAM+476 => b"00010_0011_01_0_------------", -- ADDI GR3, 13
        PROGRAM+477 => b"000000000000000000001101", -- 
        PROGRAM+478 => b"00001_0011_00_0_011010101010", -- ST 1700+6, GR3
        PROGRAM+479 => b"00000_0010_11_0_010111011100", -- LDN GR2, 1500
        PROGRAM+480 => b"00001_0010_00_0_011010101011", -- ST 1700+7, GR2
        PROGRAM+481 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+482 => b"00000_0010_00_0_011010101011", -- LD GR2, 1700+7
        PROGRAM+483 => b"00100_0010_01_0_------------", -- CMPI GR2, 0
        PROGRAM+484 => b"000000000000000000000000", -- 
        PROGRAM+485 => b"01100_----_00_0_001011100001", -- BEQ set_highlighted_grass
        PROGRAM+486 => b"00100_0010_01_0_------------", -- CMPI GR2, 1
        PROGRAM+487 => b"000000000000000000000001", -- 
        PROGRAM+488 => b"01100_----_00_0_001011111001", -- BEQ set_highlighted_monkey1
        PROGRAM+489 => b"00100_0010_01_0_------------", -- CMPI GR2, 5
        PROGRAM+490 => b"000000000000000000000101", -- 
        PROGRAM+491 => b"01100_----_00_0_001011111101", -- BEQ set_highlighted_monkey2
        PROGRAM+492 => b"00100_0010_01_0_------------", -- CMPI GR2, 9
        PROGRAM+493 => b"000000000000000000001001", -- 
        PROGRAM+494 => b"01100_----_00_0_001100000001", -- BEQ set_highlighted_monkey3
        PROGRAM+495 => b"00100_0010_01_0_------------", -- CMPI GR2, 13
        PROGRAM+496 => b"000000000000000000001101", -- 
        PROGRAM+497 => b"01100_----_00_0_001100000101", -- BEQ set_highlighted_monkey4
        PROGRAM+498 => b"00100_0010_01_0_------------", -- CMPI GR2, 17
        PROGRAM+499 => b"000000000000000000010001", -- 
        PROGRAM+500 => b"01100_----_00_0_001100001001", -- BEQ set_highlighted_monkey5
        PROGRAM+501 => b"00100_0010_01_0_------------", -- CMPI GR2, 21
        PROGRAM+502 => b"000000000000000000010101", -- 
        PROGRAM+503 => b"01100_----_00_0_001100001101", -- BEQ set_highlighted_monkey6
        PROGRAM+504 => b"00100_0010_01_0_------------", -- CMPI GR2, 25
        PROGRAM+505 => b"000000000000000000011001", -- 
        PROGRAM+506 => b"01100_----_00_0_001011100101", -- BEQ set_highlighted_path
        PROGRAM+507 => b"00100_0010_01_0_------------", -- CMPI GR2, 38
        PROGRAM+508 => b"000000000000000000100110", -- 
        PROGRAM+509 => b"01100_----_00_0_001011101101", -- BEQ set_highlighted_black
        PROGRAM+510 => b"00100_0010_01_0_------------", -- CMPI GR2, 45
        PROGRAM+511 => b"000000000000000000101101", -- 
        PROGRAM+512 => b"01100_----_00_0_001011110001", -- BEQ set_highlighted_reset
        PROGRAM+513 => b"00100_0010_01_0_------------", -- CMPI GR2, 47
        PROGRAM+514 => b"000000000000000000101111", -- 
        PROGRAM+515 => b"01100_----_00_0_001011110101", -- BEQ set_highlighted_quit
        PROGRAM+516 => b"00100_0010_01_0_------------", -- CMPI GR2, 50
        PROGRAM+517 => b"000000000000000000110010", -- 
        PROGRAM+518 => b"01100_----_00_0_001011101001", -- BEQ set_highlighted_continue
        PROGRAM+519 => b"00000_0010_01_0_------------", -- LDI GR2, 53
        PROGRAM+520 => b"000000000000000000110101", -- 
        PROGRAM+521 => b"00001_0010_11_0_010111011100", -- STN 1500,GR2
        PROGRAM+522 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+523 => b"00000_1111_01_1_------------", -- confirm_input_pick : LDI GR15, 0 // reset key input
        PROGRAM+524 => b"000000000000000000000000", -- 
        PROGRAM+525 => b"00000_1010_00_0_011010100111", -- LD GR10, 1700+3
        PROGRAM+526 => b"00010_1010_00_0_011010101000", -- ADD GR10, 1700+4
        PROGRAM+527 => b"01100_----_00_0_000100101010", -- BEQ read_input_end
        PROGRAM+528 => b"00000_0010_00_0_011010101011", -- LD GR2, 1700+7
        PROGRAM+529 => b"00100_0010_01_0_------------", -- CMPI GR2, 1
        PROGRAM+530 => b"000000000000000000000001", -- 
        PROGRAM+531 => b"00000_1001_01_0_------------", -- LDI GR9, 39
        PROGRAM+532 => b"000000000000000000100111", -- 
        PROGRAM+533 => b"01100_----_00_0_001000111011", -- BEQ confirm_input_place
        PROGRAM+534 => b"00100_0010_01_0_------------", -- CMPI GR2, 5
        PROGRAM+535 => b"000000000000000000000101", -- 
        PROGRAM+536 => b"00000_1001_01_0_------------", -- LDI GR9, 40
        PROGRAM+537 => b"000000000000000000101000", -- 
        PROGRAM+538 => b"01100_----_00_0_001000111011", -- BEQ confirm_input_place
        PROGRAM+539 => b"00100_0010_01_0_------------", -- CMPI GR2, 9
        PROGRAM+540 => b"000000000000000000001001", -- 
        PROGRAM+541 => b"00000_1001_01_0_------------", -- LDI GR9, 41
        PROGRAM+542 => b"000000000000000000101001", -- 
        PROGRAM+543 => b"01100_----_00_0_001000111011", -- BEQ confirm_input_place
        PROGRAM+544 => b"00100_0010_01_0_------------", -- CMPI GR2, 13
        PROGRAM+545 => b"000000000000000000001101", -- 
        PROGRAM+546 => b"00000_1001_01_0_------------", -- LDI GR9, 42
        PROGRAM+547 => b"000000000000000000101010", -- 
        PROGRAM+548 => b"01100_----_00_0_001000111011", -- BEQ confirm_input_place
        PROGRAM+549 => b"00100_0010_01_0_------------", -- CMPI GR2, 17
        PROGRAM+550 => b"000000000000000000010001", -- 
        PROGRAM+551 => b"00000_1001_01_0_------------", -- LDI GR9, 43
        PROGRAM+552 => b"000000000000000000101011", -- 
        PROGRAM+553 => b"01100_----_00_0_001000111011", -- BEQ confirm_input_place
        PROGRAM+554 => b"00100_0010_01_0_------------", -- CMPI GR2, 21
        PROGRAM+555 => b"000000000000000000010101", -- 
        PROGRAM+556 => b"00000_1001_01_0_------------", -- LDI GR9, 44
        PROGRAM+557 => b"000000000000000000101100", -- 
        PROGRAM+558 => b"01100_----_00_0_001000111011", -- BEQ confirm_input_place
        PROGRAM+559 => b"00000_1001_01_0_------------", -- LDI GR9, 0
        PROGRAM+560 => b"000000000000000000000000", -- 
        PROGRAM+561 => b"00100_0010_01_0_------------", -- CMPI GR2, 45 // reset
        PROGRAM+562 => b"000000000000000000101101", -- 
        PROGRAM+563 => b"01100_----_00_0_000011110001", -- BEQ dead
        PROGRAM+564 => b"00100_0010_01_0_------------", -- CMPI GR2, 47 // quit
        PROGRAM+565 => b"000000000000000000101111", -- 
        PROGRAM+566 => b"01100_----_00_0_000011110001", -- BEQ dead
        PROGRAM+567 => b"00100_0010_01_0_------------", -- CMPI GR2, 50 // continue
        PROGRAM+568 => b"000000000000000000110010", -- 
        PROGRAM+569 => b"01100_----_00_0_001010101110", -- BEQ continue_game
        PROGRAM+570 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+571 => b"01001_----_00_0_000011110010", -- confirm_input_place : JSR wait_for_break
        PROGRAM+572 => b"01001_----_00_0_000011110110", -- JSR wait_until_break_is_gone
        PROGRAM+573 => b"00100_1111_01_1_------------", -- CMPI GR15, 3 // Space
        PROGRAM+574 => b"000000000000000000000011", -- 
        PROGRAM+575 => b"01100_----_00_0_001001001101", -- BEQ place_check
        PROGRAM+576 => b"00100_1111_01_1_------------", -- CMPI GR15, 4 // W
        PROGRAM+577 => b"000000000000000000000100", -- 
        PROGRAM+578 => b"01100_----_00_0_001001111010", -- BEQ place_up
        PROGRAM+579 => b"00100_1111_01_1_------------", -- CMPI GR15, 1 // A
        PROGRAM+580 => b"000000000000000000000001", -- 
        PROGRAM+581 => b"01100_----_00_0_001010000111", -- BEQ place_left
        PROGRAM+582 => b"00100_1111_01_1_------------", -- CMPI GR15, 2 // S
        PROGRAM+583 => b"000000000000000000000010", -- 
        PROGRAM+584 => b"01100_----_00_0_001010010100", -- BEQ place_right
        PROGRAM+585 => b"00100_1111_01_1_------------", -- CMPI GR15, 8 // D
        PROGRAM+586 => b"000000000000000000001000", -- 
        PROGRAM+587 => b"01100_----_00_0_001010100001", -- BEQ place_down
        PROGRAM+588 => b"01010_----_00_0_001000111011", -- BRA confirm_input_place // Check again
        PROGRAM+589 => b"00000_0011_00_0_011010101010", -- place_check : LD GR3, 1700+6
        PROGRAM+590 => b"00000_0010_00_0_011010101011", -- LD GR2, 1700+7
        PROGRAM+591 => b"00100_0010_01_0_------------", -- CMPI GR2, 0
        PROGRAM+592 => b"000000000000000000000000", -- 
        PROGRAM+593 => b"01011_----_00_0_001000111011", -- BNE confirm_input_place // if not being placed on grass keep checking for inputs
        PROGRAM+594 => b"00100_1001_01_0_------------", -- CMPI GR9, 39
        PROGRAM+595 => b"000000000000000000100111", -- 
        PROGRAM+596 => b"00000_0010_01_0_------------", -- LDI GR2, 1
        PROGRAM+597 => b"000000000000000000000001", -- 
        PROGRAM+598 => b"01100_----_00_0_001001101101", -- BEQ purchase
        PROGRAM+599 => b"00100_1001_01_0_------------", -- CMPI GR9, 40
        PROGRAM+600 => b"000000000000000000101000", -- 
        PROGRAM+601 => b"00000_0010_01_0_------------", -- LDI GR2, 5
        PROGRAM+602 => b"000000000000000000000101", -- 
        PROGRAM+603 => b"01100_----_00_0_001001101101", -- BEQ purchase
        PROGRAM+604 => b"00100_1001_01_0_------------", -- CMPI GR9, 41
        PROGRAM+605 => b"000000000000000000101001", -- 
        PROGRAM+606 => b"00000_0010_01_0_------------", -- LDI GR2, 9
        PROGRAM+607 => b"000000000000000000001001", -- 
        PROGRAM+608 => b"01100_----_00_0_001001101101", -- BEQ purchase
        PROGRAM+609 => b"00100_1001_01_0_------------", -- CMPI GR9, 42
        PROGRAM+610 => b"000000000000000000101010", -- 
        PROGRAM+611 => b"00000_0010_01_0_------------", -- LDI GR2, 13
        PROGRAM+612 => b"000000000000000000001101", -- 
        PROGRAM+613 => b"01100_----_00_0_001001101101", -- BEQ purchase
        PROGRAM+614 => b"00100_1001_01_0_------------", -- CMPI GR9, 43
        PROGRAM+615 => b"000000000000000000101011", -- 
        PROGRAM+616 => b"00000_0010_01_0_------------", -- LDI GR2, 17
        PROGRAM+617 => b"000000000000000000010001", -- 
        PROGRAM+618 => b"01100_----_00_0_001001101101", -- BEQ purchase
        PROGRAM+619 => b"00000_0010_01_0_------------", -- LDI GR2, 21
        PROGRAM+620 => b"000000000000000000010101", -- 
        PROGRAM+621 => b"00000_1010_00_0_011010100111", -- purchase : LD GR10, 1700+3
        PROGRAM+622 => b"00100_1010_01_0_------------", -- CMPI GR10, 0
        PROGRAM+623 => b"000000000000000000000000", -- 
        PROGRAM+624 => b"01100_----_00_0_001010111100", -- BEQ decrement_of_gold
        PROGRAM+625 => b"00011_1010_01_0_------------", -- SUBI GR10, 1
        PROGRAM+626 => b"000000000000000000000001", -- 
        PROGRAM+627 => b"00001_1010_00_0_011010100111", -- ST 1700+3, GR10
        PROGRAM+628 => b"01001_----_00_0_000100111000", -- place : JSR update_gold
        PROGRAM+629 => b"00001_0010_00_0_011010101011", -- ST 1700+7, GR2
        PROGRAM+630 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+631 => b"00000_1111_01_1_------------", -- LDI GR15, 0
        PROGRAM+632 => b"000000000000000000000000", -- 
        PROGRAM+633 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+634 => b"00000_0010_00_0_011010101011", -- place_up : LD GR2, 1700+7
        PROGRAM+635 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+636 => b"00001_0010_11_0_010111011100", -- STN 1500,GR2
        PROGRAM+637 => b"00011_0011_01_0_------------", -- SUBI GR3, 13
        PROGRAM+638 => b"000000000000000000001101", -- 
        PROGRAM+639 => b"00001_0011_00_0_011010101010", -- ST 1700+6, GR3
        PROGRAM+640 => b"00000_0010_11_0_010111011100", -- LDN GR2, 1500
        PROGRAM+641 => b"00001_0010_00_0_011010101011", -- ST 1700+7, GR2
        PROGRAM+642 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+643 => b"00001_1001_11_0_010111011100", -- STN 1500, GR9
        PROGRAM+644 => b"00000_1111_01_1_------------", -- LDI GR15, 0
        PROGRAM+645 => b"000000000000000000000000", -- 
        PROGRAM+646 => b"01010_----_00_0_001000111011", -- BRA confirm_input_place
        PROGRAM+647 => b"00000_0010_00_0_011010101011", -- place_left : LD GR2, 1700+7
        PROGRAM+648 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+649 => b"00001_0010_11_0_010111011100", -- STN 1500,GR2
        PROGRAM+650 => b"00011_0011_01_0_------------", -- SUBI GR3, 1
        PROGRAM+651 => b"000000000000000000000001", -- 
        PROGRAM+652 => b"00001_0011_00_0_011010101010", -- ST 1700+6, GR3
        PROGRAM+653 => b"00000_0010_11_0_010111011100", -- LDN GR2, 1500
        PROGRAM+654 => b"00001_0010_00_0_011010101011", -- ST 1700+7, GR2
        PROGRAM+655 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+656 => b"00001_1001_11_0_010111011100", -- STN 1500, GR9
        PROGRAM+657 => b"00000_1111_01_1_------------", -- LDI GR15, 0
        PROGRAM+658 => b"000000000000000000000000", -- 
        PROGRAM+659 => b"01010_----_00_0_001000111011", -- BRA confirm_input_place
        PROGRAM+660 => b"00000_0010_00_0_011010101011", -- place_right : LD GR2, 1700+7
        PROGRAM+661 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+662 => b"00001_0010_11_0_010111011100", -- STN 1500,GR2
        PROGRAM+663 => b"00010_0011_01_0_------------", -- ADDI GR3, 1
        PROGRAM+664 => b"000000000000000000000001", -- 
        PROGRAM+665 => b"00001_0011_00_0_011010101010", -- ST 1700+6, GR3
        PROGRAM+666 => b"00000_0010_11_0_010111011100", -- LDN GR2, 1500
        PROGRAM+667 => b"00001_0010_00_0_011010101011", -- ST 1700+7, GR2
        PROGRAM+668 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+669 => b"00001_1001_11_0_010111011100", -- STN 1500, GR9
        PROGRAM+670 => b"00000_1111_01_1_------------", -- LDI GR15, 0
        PROGRAM+671 => b"000000000000000000000000", -- 
        PROGRAM+672 => b"01010_----_00_0_001000111011", -- BRA confirm_input_place
        PROGRAM+673 => b"00000_0010_00_0_011010101011", -- place_down : LD GR2, 1700+7
        PROGRAM+674 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+675 => b"00001_0010_11_0_010111011100", -- STN 1500,GR2
        PROGRAM+676 => b"00010_0011_01_0_------------", -- ADDI GR3, 13
        PROGRAM+677 => b"000000000000000000001101", -- 
        PROGRAM+678 => b"00001_0011_00_0_011010101010", -- ST 1700+6, GR3
        PROGRAM+679 => b"00000_0010_11_0_010111011100", -- LDN GR2, 1500
        PROGRAM+680 => b"00001_0010_00_0_011010101011", -- ST 1700+7, GR2
        PROGRAM+681 => b"00000_0011_00_0_011010101010", -- LD GR3, 1700+6
        PROGRAM+682 => b"00001_1001_11_0_010111011100", -- STN 1500, GR9
        PROGRAM+683 => b"00000_1111_01_1_------------", -- LDI GR15, 0
        PROGRAM+684 => b"000000000000000000000000", -- 
        PROGRAM+685 => b"01010_----_00_0_001000111011", -- BRA confirm_input_place
        PROGRAM+686 => b"00000_0011_00_0_011010101010", -- continue_game : LD GR3, 1700+6
        PROGRAM+687 => b"00000_0010_00_0_011010101011", -- LD GR2, 1700+7
        PROGRAM+688 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+689 => b"00000_1000_01_0_------------", -- LDI GR8, 1
        PROGRAM+690 => b"000000000000000000000001", -- 
        PROGRAM+691 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+692 => b"00000_0111_01_0_------------", -- increment_of_gold : LDI GR7, 0
        PROGRAM+693 => b"000000000000000000000000", -- 
        PROGRAM+694 => b"00001_0111_00_0_011010100111", -- ST 1700+3, GR7
        PROGRAM+695 => b"00000_0111_00_0_011010101000", -- LD GR7, 1700+4
        PROGRAM+696 => b"00010_0111_01_0_------------", -- ADDI GR7, 1
        PROGRAM+697 => b"000000000000000000000001", -- 
        PROGRAM+698 => b"00001_0111_00_0_011010101000", -- ST 1700+4, GR7
        PROGRAM+699 => b"01010_----_00_0_000010111110", -- BRA balloon_dead2
        PROGRAM+700 => b"00000_0111_00_0_011010101000", -- decrement_of_gold : LD GR7, 1700+4
        PROGRAM+701 => b"00100_0111_01_0_------------", -- CMPI GR7, 0
        PROGRAM+702 => b"000000000000000000000000", -- 
        PROGRAM+703 => b"01100_----_00_0_001000111011", -- BEQ confirm_input_place
        PROGRAM+704 => b"00000_1010_01_0_------------", -- LDI GR10, 9
        PROGRAM+705 => b"000000000000000000001001", -- 
        PROGRAM+706 => b"00001_1010_00_0_011010100111", -- ST 1700+3, GR10
        PROGRAM+707 => b"00000_1010_00_0_011010101000", -- LD GR10, 1700+4
        PROGRAM+708 => b"00011_1010_01_0_------------", -- SUBI GR10, 1
        PROGRAM+709 => b"000000000000000000000001", -- 
        PROGRAM+710 => b"00001_1010_00_0_011010101000", -- ST 1700+4, GR10
        PROGRAM+711 => b"01010_----_00_0_001001110100", -- BRA place
        PROGRAM+712 => b"00000_0111_00_0_011010100110", -- decrement_of_hp : LD GR7, 1700+2
        PROGRAM+713 => b"00100_0111_01_0_------------", -- CMPI GR7, 0
        PROGRAM+714 => b"000000000000000000000000", -- 
        PROGRAM+715 => b"01100_----_00_0_000010100001", -- BEQ player_dmg_2
        PROGRAM+716 => b"00000_0010_01_0_------------", -- LDI GR2, 9
        PROGRAM+717 => b"000000000000000000001001", -- 
        PROGRAM+718 => b"00001_0010_00_0_011010100101", -- ST 1700+1, GR2
        PROGRAM+719 => b"00000_0010_00_0_011010100110", -- LD GR2, 1700+2
        PROGRAM+720 => b"00011_0010_01_0_------------", -- SUBI GR2, 1
        PROGRAM+721 => b"000000000000000000000001", -- 
        PROGRAM+722 => b"00001_0010_00_0_011010100110", -- ST 1700+2, GR2
        PROGRAM+723 => b"01010_----_00_0_000010100001", -- BRA player_dmg_2
        PROGRAM+724 => b"01101_0000_--_0_------------", -- delay : PUSH GR0
        PROGRAM+725 => b"00000_0000_00_0_011010101100", -- LD GR0, 1700+8
        PROGRAM+726 => b"00011_0000_01_0_------------", -- delay_loop : SUBI GR0, 1
        PROGRAM+727 => b"000000000000000000000001", -- 
        PROGRAM+728 => b"01011_----_00_0_001011010110", -- BNE delay_loop
        PROGRAM+729 => b"01110_0000_--_0_------------", -- delay_end : POP GR0
        PROGRAM+730 => b"10000_----_--_0_------------", -- RET
        PROGRAM+731 => b"00100_1111_01_1_------------", -- wait_for_player_input : CMPI GR15, 3     // loop until user input
        PROGRAM+732 => b"000000000000000000000011", -- 
        PROGRAM+733 => b"01011_----_00_0_001011011011", -- BNE wait_for_player_input
        PROGRAM+734 => b"00000_1111_01_1_------------", -- LDI GR15, 0
        PROGRAM+735 => b"000000000000000000000000", -- 
        PROGRAM+736 => b"10000_----_--_0_------------", -- RET
        PROGRAM+737 => b"00000_0010_01_0_------------", -- set_highlighted_grass : LDI GR2, 65
        PROGRAM+738 => b"000000000000000001000001", -- 
        PROGRAM+739 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+740 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+741 => b"00000_0010_01_0_------------", -- set_highlighted_path : LDI GR2, 66
        PROGRAM+742 => b"000000000000000001000010", -- 
        PROGRAM+743 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+744 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+745 => b"00000_0010_01_0_------------", -- set_highlighted_continue : LDI GR2, 52
        PROGRAM+746 => b"000000000000000000110100", -- 
        PROGRAM+747 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+748 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+749 => b"00000_0010_01_0_------------", -- set_highlighted_black : LDI GR2, 53
        PROGRAM+750 => b"000000000000000000110101", -- 
        PROGRAM+751 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+752 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+753 => b"00000_0010_01_0_------------", -- set_highlighted_reset : LDI GR2, 46
        PROGRAM+754 => b"000000000000000000101110", -- 
        PROGRAM+755 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+756 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+757 => b"00000_0010_01_0_------------", -- set_highlighted_quit : LDI GR2, 48
        PROGRAM+758 => b"000000000000000000110000", -- 
        PROGRAM+759 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+760 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+761 => b"00000_0010_01_0_------------", -- set_highlighted_monkey1 : LDI GR2, 39
        PROGRAM+762 => b"000000000000000000100111", -- 
        PROGRAM+763 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+764 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+765 => b"00000_0010_01_0_------------", -- set_highlighted_monkey2 : LDI GR2, 40
        PROGRAM+766 => b"000000000000000000101000", -- 
        PROGRAM+767 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+768 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+769 => b"00000_0010_01_0_------------", -- set_highlighted_monkey3 : LDI GR2, 41
        PROGRAM+770 => b"000000000000000000101001", -- 
        PROGRAM+771 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+772 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+773 => b"00000_0010_01_0_------------", -- set_highlighted_monkey4 : LDI GR2, 42
        PROGRAM+774 => b"000000000000000000101010", -- 
        PROGRAM+775 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+776 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+777 => b"00000_0010_01_0_------------", -- set_highlighted_monkey5 : LDI GR2, 43
        PROGRAM+778 => b"000000000000000000101011", -- 
        PROGRAM+779 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+780 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        PROGRAM+781 => b"00000_0010_01_0_------------", -- set_highlighted_monkey6 : LDI GR2, 44
        PROGRAM+782 => b"000000000000000000101100", -- 
        PROGRAM+783 => b"00001_0010_11_0_010111011100", -- STN 1500, GR2
        PROGRAM+784 => b"01010_----_00_0_000100101010", -- BRA read_input_end
        -- VMEM
        VMEM+0 => b"000000000000000000000000", -- 0
        VMEM+1 => b"000000000000000000000000", -- 0
        VMEM+2 => b"000000000000000000000000", -- 0
        VMEM+3 => b"000000000000000000000000", -- 0
        VMEM+4 => b"000000000000000000000000", -- 0
        VMEM+5 => b"000000000000000000000000", -- 0
        VMEM+6 => b"000000000000000000000000", -- 0
        VMEM+7 => b"000000000000000000000000", -- 0
        VMEM+8 => b"000000000000000000000000", -- 0
        VMEM+9 => b"000000000000000000000000", -- 0
        VMEM+10 => b"000000000000000000110001", -- 49
        VMEM+11 => b"000000000000000000111111", -- 63
        VMEM+12 => b"000000000000000000111111", -- 63
        VMEM+13 => b"000000000000000000000000", -- 0
        VMEM+14 => b"000000000000000000011001", -- 25
        VMEM+15 => b"000000000000000000011001", -- 25
        VMEM+16 => b"000000000000000000011001", -- 25
        VMEM+17 => b"000000000000000000011001", -- 25
        VMEM+18 => b"000000000000000000011001", -- 25
        VMEM+19 => b"000000000000000000011001", -- 25
        VMEM+20 => b"000000000000000000011001", -- 25
        VMEM+21 => b"000000000000000000011001", -- 25
        VMEM+22 => b"000000000000000000000000", -- 0
        VMEM+23 => b"000000000000000000110011", -- 51
        VMEM+24 => b"000000000000000000110110", -- 54
        VMEM+25 => b"000000000000000000110110", -- 54
        VMEM+26 => b"000000000000000000000000", -- 0
        VMEM+27 => b"000000000000000000011001", -- 25
        VMEM+28 => b"000000000000000000000000", -- 0
        VMEM+29 => b"000000000000000000000000", -- 0
        VMEM+30 => b"000000000000000000000000", -- 0
        VMEM+31 => b"000000000000000000000000", -- 0
        VMEM+32 => b"000000000000000000000000", -- 0
        VMEM+33 => b"000000000000000000000000", -- 0
        VMEM+34 => b"000000000000000000011001", -- 25
        VMEM+35 => b"000000000000000000000000", -- 0
        VMEM+36 => b"000000000000000000000001", -- 1
        VMEM+37 => b"000000000000000000100110", -- 38
        VMEM+38 => b"000000000000000000000101", -- 5
        VMEM+39 => b"000000000000000000000000", -- 0
        VMEM+40 => b"000000000000000000011001", -- 25
        VMEM+41 => b"000000000000000000000000", -- 0
        VMEM+42 => b"000000000000000000011001", -- 25
        VMEM+43 => b"000000000000000000011001", -- 25
        VMEM+44 => b"000000000000000000011001", -- 25
        VMEM+45 => b"000000000000000000011001", -- 25
        VMEM+46 => b"000000000000000000011001", -- 25
        VMEM+47 => b"000000000000000000011001", -- 25
        VMEM+48 => b"000000000000000000000000", -- 0
        VMEM+49 => b"000000000000000000100110", -- 38
        VMEM+50 => b"000000000000000000100110", -- 38
        VMEM+51 => b"000000000000000000100110", -- 38
        VMEM+52 => b"000000000000000000011001", -- 25
        VMEM+53 => b"000000000000000000011001", -- 25
        VMEM+54 => b"000000000000000000000000", -- 0
        VMEM+55 => b"000000000000000000011001", -- 25
        VMEM+56 => b"000000000000000000000000", -- 0
        VMEM+57 => b"000000000000000000000000", -- 0
        VMEM+58 => b"000000000000000000000000", -- 0
        VMEM+59 => b"000000000000000000000000", -- 0
        VMEM+60 => b"000000000000000000000000", -- 0
        VMEM+61 => b"000000000000000000000000", -- 0
        VMEM+62 => b"000000000000000000001001", -- 9
        VMEM+63 => b"000000000000000000100110", -- 38
        VMEM+64 => b"000000000000000000001101", -- 13
        VMEM+65 => b"000000000000000000000000", -- 0
        VMEM+66 => b"000000000000000000000000", -- 0
        VMEM+67 => b"000000000000000000000000", -- 0
        VMEM+68 => b"000000000000000000011001", -- 25
        VMEM+69 => b"000000000000000000000000", -- 0
        VMEM+70 => b"000000000000000000011001", -- 25
        VMEM+71 => b"000000000000000000011001", -- 25
        VMEM+72 => b"000000000000000000011001", -- 25
        VMEM+73 => b"000000000000000000000000", -- 0
        VMEM+74 => b"000000000000000000000000", -- 0
        VMEM+75 => b"000000000000000000100110", -- 38
        VMEM+76 => b"000000000000000000100110", -- 38
        VMEM+77 => b"000000000000000000100110", -- 38
        VMEM+78 => b"000000000000000000000000", -- 0
        VMEM+79 => b"000000000000000000011001", -- 25
        VMEM+80 => b"000000000000000000011001", -- 25
        VMEM+81 => b"000000000000000000011001", -- 25
        VMEM+82 => b"000000000000000000000000", -- 0
        VMEM+83 => b"000000000000000000011001", -- 25
        VMEM+84 => b"000000000000000000000000", -- 0
        VMEM+85 => b"000000000000000000011001", -- 25
        VMEM+86 => b"000000000000000000000000", -- 0
        VMEM+87 => b"000000000000000000000000", -- 0
        VMEM+88 => b"000000000000000000010001", -- 17
        VMEM+89 => b"000000000000000000100110", -- 38
        VMEM+90 => b"000000000000000000010101", -- 21
        VMEM+91 => b"000000000000000000000000", -- 0
        VMEM+92 => b"000000000000000000011001", -- 25
        VMEM+93 => b"000000000000000000000000", -- 0
        VMEM+94 => b"000000000000000000000000", -- 0
        VMEM+95 => b"000000000000000000000000", -- 0
        VMEM+96 => b"000000000000000000011001", -- 25
        VMEM+97 => b"000000000000000000000000", -- 0
        VMEM+98 => b"000000000000000000011001", -- 25
        VMEM+99 => b"000000000000000000000000", -- 0
        VMEM+100 => b"000000000000000000000000", -- 0
        VMEM+101 => b"000000000000000000100110", -- 38
        VMEM+102 => b"000000000000000000100110", -- 38
        VMEM+103 => b"000000000000000000100110", -- 38
        VMEM+104 => b"000000000000000000000000", -- 0
        VMEM+105 => b"000000000000000000011001", -- 25
        VMEM+106 => b"000000000000000000011001", -- 25
        VMEM+107 => b"000000000000000000011001", -- 25
        VMEM+108 => b"000000000000000000011001", -- 25
        VMEM+109 => b"000000000000000000011001", -- 25
        VMEM+110 => b"000000000000000000000000", -- 0
        VMEM+111 => b"000000000000000000011001", -- 25
        VMEM+112 => b"000000000000000000011001", -- 25
        VMEM+113 => b"000000000000000000011001", -- 25
        VMEM+114 => b"000000000000000000100110", -- 38
        VMEM+115 => b"000000000000000000100110", -- 38
        VMEM+116 => b"000000000000000000100110", -- 38
        VMEM+117 => b"000000000000000000000000", -- 0
        VMEM+118 => b"000000000000000000000000", -- 0
        VMEM+119 => b"000000000000000000000000", -- 0
        VMEM+120 => b"000000000000000000000000", -- 0
        VMEM+121 => b"000000000000000000000000", -- 0
        VMEM+122 => b"000000000000000000000000", -- 0
        VMEM+123 => b"000000000000000000000000", -- 0
        VMEM+124 => b"000000000000000000000000", -- 0
        VMEM+125 => b"000000000000000000000000", -- 0
        VMEM+126 => b"000000000000000000000000", -- 0
        VMEM+127 => b"000000000000000000101101", -- 45
        VMEM+128 => b"000000000000000000110010", -- 50
        VMEM+129 => b"000000000000000000101111", -- 47
        -- PATH
        PATH+0 => b"000000000000000000110100", -- 52
        PATH+1 => b"000000000000000000110101", -- 53
        PATH+2 => b"000000000000000000101000", -- 40
        PATH+3 => b"000000000000000000011011", -- 27
        PATH+4 => b"000000000000000000001110", -- 14
        PATH+5 => b"000000000000000000001111", -- 15
        PATH+6 => b"000000000000000000010000", -- 16
        PATH+7 => b"000000000000000000010001", -- 17
        PATH+8 => b"000000000000000000010010", -- 18
        PATH+9 => b"000000000000000000010011", -- 19
        PATH+10 => b"000000000000000000010100", -- 20
        PATH+11 => b"000000000000000000010101", -- 21
        PATH+12 => b"000000000000000000100010", -- 34
        PATH+13 => b"000000000000000000101111", -- 47
        PATH+14 => b"000000000000000000101110", -- 46
        PATH+15 => b"000000000000000000101101", -- 45
        PATH+16 => b"000000000000000000101100", -- 44
        PATH+17 => b"000000000000000000101011", -- 43
        PATH+18 => b"000000000000000000101010", -- 42
        PATH+19 => b"000000000000000000110111", -- 55
        PATH+20 => b"000000000000000001000100", -- 68
        PATH+21 => b"000000000000000001010001", -- 81
        PATH+22 => b"000000000000000001010000", -- 80
        PATH+23 => b"000000000000000001001111", -- 79
        PATH+24 => b"000000000000000001011100", -- 92
        PATH+25 => b"000000000000000001101001", -- 105
        PATH+26 => b"000000000000000001101010", -- 106
        PATH+27 => b"000000000000000001101011", -- 107
        PATH+28 => b"000000000000000001101100", -- 108
        PATH+29 => b"000000000000000001101101", -- 109
        PATH+30 => b"000000000000000001100000", -- 96
        PATH+31 => b"000000000000000001010011", -- 83
        PATH+32 => b"000000000000000001000110", -- 70
        PATH+33 => b"000000000000000001000111", -- 71
        PATH+34 => b"000000000000000001001000", -- 72
        PATH+35 => b"000000000000000001010101", -- 85
        PATH+36 => b"000000000000000001100010", -- 98
        PATH+37 => b"000000000000000001101111", -- 111
        PATH+38 => b"000000000000000001110000", -- 112
        PATH+39 => b"000000000000000001110001", -- 113
        PATH+40 => b"000000000000000001110010", -- 114
        -- HEAP
        OTHERS => (OTHERS => '-')
    );

BEGIN

    -- Reading from two-port ram
    PROCESS (clk)
    BEGIN
        IF rising_edge(clk) THEN
            cpu_data_out <= p_mem(TO_INTEGER(cpu_address) + PROGRAM);
            video_data_out <= unsigned(p_mem(TO_INTEGER(video_address) + VMEM)(6 DOWNTO 0));
        END IF;
    END PROCESS;

    -- STORE
    PROCESS (clk)
    BEGIN
        IF rising_edge(clk) THEN
            IF (cpu_we = '1') THEN
                p_mem(TO_INTEGER(cpu_address)) <= STD_LOGIC_VECTOR(cpu_data_in);
            END IF;
        END IF;
    END PROCESS;

END ARCHITECTURE;