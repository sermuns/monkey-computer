LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY tile_rom IS
    PORT (
        address : IN UNSIGNED(13 DOWNTO 0); -- 14 bit address
        data_out : OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
    );
END tile_rom;

ARCHITECTURE func OF tile_rom IS
    TYPE palette_rom_type IS ARRAY(0 TO 31) OF STD_LOGIC_VECTOR(11 DOWNTO 0);
    CONSTANT palette_rom : palette_rom_type := (
        00 => x"fff",
        01 => x"000",
        02 => x"322",
        03 => x"444",
        04 => x"fa9",
        05 => x"743",
        06 => x"931",
        07 => x"c85",
        08 => x"fd5",
        09 => x"160",
        10 => x"4eb",
        11 => x"38d",
        12 => x"000",
        13 => x"557",
        14 => x"54a",
        15 => x"423",
        16 => x"712",
        17 => x"e67",
        18 => x"b22",
        19 => x"UUU",
        20 => x"UUU",
        21 => x"UUU",
        22 => x"UUU",
        23 => x"UUU",
        24 => x"UUU",
        25 => x"UUU",
        26 => x"UUU",
        27 => x"UUU",
        28 => x"UUU",
        29 => x"UUU",
        30 => x"UUU",
        31 => x"UUU"
    );

    CONSTANT NUM_TILES : INTEGER := 32;
    CONSTANT TILE_SIZE : INTEGER := 12*12;

    TYPE tile_rom_type IS ARRAY(0 TO TILE_SIZE*NUM_TILES) OF unsigned(4 DOWNTO 0);
    CONSTANT tile_rom_data : tile_rom_type := (
        -- 0
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00000",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "01110", "01011", "00000", "00000", "01110", "01011", "00000", "00000", "00000",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        -- 1
        "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00000",
        "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00000",
        "00001", "00001", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00111", "00111", "00000", "00000", "00111", "00111", "00000", "00000", "00000",
        "00000", "00000", "00000", "00111", "00111", "00000", "00000", "00111", "00111", "00000", "00000", "00000",
        "00000", "00000", "00000", "00111", "00111", "00000", "00000", "00111", "00111", "00000", "00000", "00000",
        "00000", "00000", "00000", "00111", "00111", "00000", "00000", "00111", "00111", "00000", "00000", "00000",
        "00000", "00000", "01011", "00110", "00110", "01110", "01011", "00110", "00110", "01110", "00000", "00000",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "00000", "00000", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00000", "00000",
        "00000", "00001", "00000", "00101", "00101", "00000", "00000", "00101", "00101", "00000", "00000", "00000",
        -- 2
        "00001", "00001", "00000", "00101", "00101", "00000", "00000", "00101", "00101", "00000", "00000", "00000",
        "00000", "00000", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "00000", "00000",
        "00000", "00000", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "00000", "00000",
        "00000", "00000", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "00000", "00000",
        "00000", "00000", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "00000", "00000",
        "00000", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "00000",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "00000", "00000", "00101", "00101", "00001", "00101", "00101", "00001", "00101", "00101", "00000", "00000",
        "00000", "00000", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00000", "00000",
        "00000", "00000", "00000", "00101", "00101", "00000", "00000", "00101", "00101", "00000", "00000", "00000",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00000", "00000",

        OTHERS => (OTHERS => 'U')
    );

    SIGNAL palette_index : unsigned(4 DOWNTO 0); -- max 32 colors
BEGIN
    PROCESS (address)
    BEGIN
        -- get palette index from memory
        palette_index <= tile_rom_data(to_integer(address));
        data_out <= palette_rom(to_integer(palette_index));
    END PROCESS;
END ARCHITECTURE;