LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

-- usage: 
-- give uAddr, get uData at that address
ENTITY uMem IS
    PORT (
        uAddr : IN unsigned(7 DOWNTO 0);
        uData : OUT unsigned(23 DOWNTO 0));
END uMem;

ARCHITECTURE func OF uMem IS
    TYPE u_mem_t IS ARRAY(1000 DOWNTO 0) OF unsigned(23 DOWNTO 0);
    CONSTANT u_mem_c : u_mem_t :=
    -- "000_000_0000_0_0000_000000000" = "TB_FB_ALU_P_SEQ_uADR"
    (
    b"010_000_0000_0_0000_000000000", -- ASR := PC
    b"001_100_0000_1_0101_000000000", -- IR := PM, PC := PC + 1, uPC := uADR  
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000",
    b"000_000_0000_0_0000_000000000"
    );
    SIGNAL u_mem : u_mem_t := u_mem_c;

BEGIN
    uData <= u_mem(TO_INTEGER(uAddr));
END ARCHITECTURE;