LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY tile_rom IS
    PORT (
        clk : IN STD_LOGIC;
        address : IN UNSIGNED(13 DOWNTO 0); -- 14 bit address
        data_out : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
    );
END tile_rom;

ARCHITECTURE func OF tile_rom IS TYPE palette_rom_type IS ARRAY(0 TO 18) OF STD_LOGIC_VECTOR(23 DOWNTO 0);
    CONSTANT palette_rom : palette_rom_type := (
        00 => x"000000",
        01 => x"ffffff",
        02 => x"332222",
        03 => x"404040",
        04 => x"f5a097",
        05 => x"774433",
        06 => x"993311",
        07 => x"cc8855",
        08 => x"ffdd55",
        09 => x"176b04",
        10 => x"44eebb",
        11 => x"3388dd",
        12 => x"070708",
        13 => x"555577",
        14 => x"5544aa",
        15 => x"422433",
        16 => x"73172d",
        17 => x"e86a73",
        18 => x"b4202a"
    );
    CONSTANT TILE_SIZE : INTEGER := 12 * 12;

    TYPE tile_rom_type IS ARRAY(0 TO 7487) OF unsigned(4 DOWNTO 0);
    CONSTANT tile_rom_data : tile_rom_type := (
        -- 0
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        -- 1
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00000", "00000", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00001", "00101", "00101", "00101", "00101", "00001", "00101", "00001", "00001",
        "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        -- 2
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00000", "00000", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00001", "00101", "00101", "00101", "00101", "00001", "00101", "00001", "00001",
        "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        -- 3
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00000", "00000", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00001", "00101", "00101", "00101", "00101", "00001", "00101", "00001", "00001",
        "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        -- 4
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00000", "00000", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00001", "00101", "00101", "00101", "00101", "00001", "00101", "00001", "00001",
        "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        -- 5
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00111", "00111", "00001", "00001", "00111", "00111", "00001", "00001", "00001",
        "00001", "00001", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "00001", "00001",
        "00001", "00001", "00111", "00111", "00000", "00111", "00111", "00000", "00111", "00111", "00001", "00001",
        "00001", "00001", "00001", "00111", "00111", "00111", "00111", "00111", "00111", "00001", "01000", "00001",
        "00001", "00001", "00001", "00111", "00111", "00000", "00000", "00111", "00111", "00001", "00001", "00001",
        "00001", "00001", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00001", "00001",
        "00001", "00001", "00111", "00001", "00111", "00111", "00111", "00111", "00001", "00111", "00001", "00001",
        "00001", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00111", "00111", "00001", "00001", "00111", "00111", "00001", "00001", "00001",
        -- 6
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00111", "00111", "00001", "00001", "00111", "00111", "00001", "00001", "00001",
        "00001", "00001", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "00001", "00001",
        "00001", "00001", "00111", "00111", "00000", "00111", "00111", "00000", "00111", "00111", "00001", "00001",
        "00001", "00001", "00001", "00111", "00111", "00111", "00111", "00111", "00111", "00001", "01000", "00001",
        "00001", "00001", "00001", "00111", "00111", "00000", "00000", "00111", "00111", "00001", "00001", "00001",
        "00001", "00001", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00001", "00001",
        "00001", "00001", "00111", "00001", "00111", "00111", "00111", "00111", "00001", "00111", "00001", "00001",
        "00001", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00111", "00001", "00001", "00001",
        "00001", "00001", "00001", "00111", "00111", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        -- 7
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00111", "00111", "00001", "00001", "00111", "00111", "00001", "00001", "00001",
        "00001", "00001", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "00001", "00001",
        "00001", "00001", "00111", "00111", "00000", "00111", "00111", "00000", "00111", "00111", "00001", "00001",
        "00001", "00001", "00001", "00111", "00111", "00111", "00111", "00111", "00111", "00001", "01000", "00001",
        "00001", "00001", "00001", "00111", "00111", "00000", "00000", "00111", "00111", "00001", "00001", "00001",
        "00001", "00001", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00001", "00001",
        "00001", "00001", "00111", "00001", "00111", "00111", "00111", "00111", "00001", "00111", "00001", "00001",
        "00001", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00111", "00111", "00001", "00001", "00111", "00111", "00001", "00001", "00001",
        -- 8
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00111", "00111", "00001", "00001", "00111", "00111", "00001", "00001", "00001",
        "00001", "00001", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "00001", "00001",
        "00001", "00001", "00111", "00111", "00000", "00111", "00111", "00000", "00111", "00111", "00001", "00001",
        "00001", "00001", "00001", "00111", "00111", "00111", "00111", "00111", "00111", "00001", "01000", "00001",
        "00001", "00001", "00001", "00111", "00111", "00000", "00000", "00111", "00111", "00001", "00001", "00001",
        "00001", "00001", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00001", "00001",
        "00001", "00001", "00111", "00001", "00111", "00111", "00111", "00111", "00001", "00111", "00001", "00001",
        "00001", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00111", "00001", "00001", "00001",
        "00001", "00001", "00001", "00111", "00111", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        -- 9
        "00001", "00001", "00001", "01110", "01011", "00001", "00001", "01110", "01011", "00001", "00001", "00001",
        "00001", "00001", "01011", "00110", "00110", "01110", "01011", "00110", "00110", "01110", "00001", "00001",
        "00001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "00001",
        "00001", "01011", "00110", "00110", "00000", "00110", "00110", "00000", "00110", "00110", "01110", "00001",
        "00001", "00001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "00001", "00001",
        "00001", "00001", "01011", "00110", "00110", "00000", "00000", "00110", "00110", "01110", "00001", "00001",
        "00001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "00001",
        "00001", "01011", "00110", "01011", "00110", "00110", "00110", "00110", "01110", "00110", "01110", "00001",
        "00001", "00001", "01110", "00001", "00110", "00001", "00001", "00110", "00001", "01011", "00001", "00001",
        "00001", "00001", "00001", "00001", "00110", "00001", "00001", "00110", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01101", "00001", "00001", "01101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "01101", "01101", "00001", "00001", "01101", "01101", "00001", "00001", "00001",
        -- 10
        "00001", "00001", "00001", "01011", "01110", "00001", "00001", "01011", "01110", "00001", "00001", "00001",
        "00001", "00001", "01110", "00110", "00110", "01011", "01110", "00110", "00110", "01011", "00001", "00001",
        "00001", "01011", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01110", "00001",
        "00001", "01110", "00110", "00110", "00000", "00110", "00110", "00000", "00110", "00110", "01011", "00001",
        "00001", "00001", "01011", "00110", "00110", "00110", "00110", "00110", "00110", "01110", "00001", "00001",
        "00001", "00001", "01110", "00110", "00110", "00000", "00000", "00110", "00110", "01011", "00001", "00001",
        "00001", "01011", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01110", "00001",
        "00001", "01110", "00110", "01110", "00110", "00110", "00110", "00110", "01011", "00110", "01011", "00001",
        "00001", "00001", "01011", "00001", "00110", "00001", "00001", "00110", "00001", "01110", "00001", "00001",
        "00001", "00001", "00001", "00001", "00110", "00001", "00001", "00110", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01101", "00001", "00001", "01101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "01101", "01101", "00001", "00001", "01101", "01101", "00001", "00001", "00001",
        -- 11
        "00001", "00001", "00001", "01110", "01011", "00001", "00001", "01110", "01011", "00001", "00001", "00001",
        "00001", "00001", "01011", "00110", "00110", "01110", "01011", "00110", "00110", "01110", "00001", "00001",
        "00001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "00001",
        "00001", "01011", "00110", "00110", "00000", "00110", "00110", "00000", "00110", "00110", "01110", "00001",
        "00001", "00001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "00001", "00001",
        "00001", "00001", "01011", "00110", "00110", "00000", "00000", "00110", "00110", "01110", "00001", "00001",
        "00001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "00001",
        "00001", "01011", "00110", "01011", "00110", "00110", "00110", "00110", "01110", "00110", "01110", "00001",
        "00001", "00001", "01110", "00001", "00110", "00001", "00001", "00110", "00001", "01011", "00001", "00001",
        "00001", "00001", "00001", "00001", "00110", "00001", "00001", "00110", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01101", "00001", "00001", "01101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "01101", "01101", "00001", "00001", "01101", "01101", "00001", "00001", "00001",
        -- 12
        "00001", "00001", "00001", "01011", "01110", "00001", "00001", "01011", "01110", "00001", "00001", "00001",
        "00001", "00001", "01110", "00110", "00110", "01011", "01110", "00110", "00110", "01011", "00001", "00001",
        "00001", "01011", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01110", "00001",
        "00001", "01110", "00110", "00110", "00000", "00110", "00110", "00000", "00110", "00110", "01011", "00001",
        "00001", "00001", "01011", "00110", "00110", "00110", "00110", "00110", "00110", "01110", "00001", "00001",
        "00001", "00001", "01110", "00110", "00110", "00000", "00000", "00110", "00110", "01011", "00001", "00001",
        "00001", "01011", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01110", "00001",
        "00001", "01110", "00110", "01110", "00110", "00110", "00110", "00110", "01011", "00110", "01011", "00001",
        "00001", "00001", "01011", "00001", "00110", "00001", "00001", "00110", "00001", "01110", "00001", "00001",
        "00001", "00001", "00001", "00001", "00110", "00001", "00001", "00110", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01101", "00001", "00001", "01101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "01101", "01101", "00001", "00001", "01101", "01101", "00001", "00001", "00001",
        -- 13
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "10000", "10001", "00001", "00001", "10001", "10000", "00001", "00001", "00001",
        "00001", "00001", "10000", "00100", "10001", "10001", "10001", "10001", "00100", "10000", "00001", "00001",
        "00001", "00001", "10001", "10001", "00000", "10001", "10001", "00000", "10001", "10001", "00001", "00001",
        "00001", "00001", "00001", "10001", "10001", "10001", "10001", "10001", "10001", "00001", "00001", "00001",
        "00001", "00001", "00001", "10001", "10001", "00000", "00000", "10001", "10001", "00001", "00001", "00001",
        "00001", "00001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "00001", "00001",
        "00001", "00001", "10001", "00001", "10001", "10001", "10001", "10001", "00001", "10001", "00001", "00001",
        "00001", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "10001", "10001", "00001", "00001", "10001", "10001", "00001", "00001", "00001",
        -- 14
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "10000", "10001", "00001", "00001", "10001", "10000", "00001", "00001", "00001",
        "00001", "00001", "10000", "00100", "10001", "10001", "10001", "10001", "00100", "10000", "00001", "00001",
        "00001", "00001", "10001", "10001", "00000", "10001", "10001", "00000", "10001", "10001", "00001", "00001",
        "00001", "00001", "00001", "10001", "10001", "10001", "10001", "10001", "10001", "00001", "00001", "00001",
        "00001", "00001", "00001", "10001", "10001", "00000", "00000", "10001", "10001", "00001", "00001", "00001",
        "00001", "00001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "00001", "00001",
        "00001", "00001", "10001", "00001", "10001", "10001", "10001", "10001", "00001", "10001", "00001", "00001",
        "00001", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "10001", "00001", "00001", "00001",
        "00001", "00001", "00001", "10001", "10001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        -- 15
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "10000", "10001", "00001", "00001", "10001", "10000", "00001", "00001", "00001",
        "00001", "00001", "10000", "00100", "10001", "10001", "10001", "10001", "00100", "10000", "00001", "00001",
        "00001", "00001", "10001", "10001", "00000", "10001", "10001", "00000", "10001", "10001", "00001", "00001",
        "00001", "00001", "00001", "10001", "10001", "10001", "10001", "10001", "10001", "00001", "00001", "00001",
        "00001", "00001", "00001", "10001", "10001", "00000", "00000", "10001", "10001", "00001", "00001", "00001",
        "00001", "00001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "00001", "00001",
        "00001", "00001", "10001", "00001", "10001", "10001", "10001", "10001", "00001", "10001", "00001", "00001",
        "00001", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "10001", "10001", "00001", "00001", "10001", "10001", "00001", "00001", "00001",
        -- 16
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "10000", "10001", "00001", "00001", "10001", "10000", "00001", "00001", "00001",
        "00001", "00001", "10000", "00100", "10001", "10001", "10001", "10001", "00100", "10000", "00001", "00001",
        "00001", "00001", "10001", "10001", "00000", "10001", "10001", "00000", "10001", "10001", "00001", "00001",
        "00001", "00001", "00001", "10001", "10001", "10001", "10001", "10001", "10001", "00001", "00001", "00001",
        "00001", "00001", "00001", "10001", "10001", "00000", "00000", "10001", "10001", "00001", "00001", "00001",
        "00001", "00001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "00001", "00001",
        "00001", "00001", "10001", "00001", "10001", "10001", "10001", "10001", "00001", "10001", "00001", "00001",
        "00001", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "10001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "10001", "10001", "00001", "00001", "00001",
        -- 17
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "00001", "00001", "01111", "01111", "00001", "00001", "00001",
        "00001", "00001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "00001", "00001",
        "00001", "00001", "01111", "01111", "00000", "01111", "01111", "00000", "01111", "01111", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "01111", "01111", "01111", "01111", "00001", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "00000", "00000", "01111", "01111", "00001", "00001", "00001",
        "00001", "00001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "00001", "00001",
        "00001", "00001", "01111", "00001", "01111", "01111", "01111", "01111", "00001", "01111", "00001", "00001",
        "00001", "00001", "00001", "00001", "01111", "00001", "00001", "01111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01111", "00001", "00001", "01111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01111", "00001", "00001", "01111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "00001", "00001", "01111", "01111", "00001", "00001", "00001",
        -- 18
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "00001", "00001", "01111", "01111", "00001", "00001", "00001",
        "00001", "00001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "00001", "00001",
        "00001", "00001", "01111", "01111", "00000", "01111", "01111", "00000", "01111", "01111", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "01111", "01111", "01111", "01111", "00001", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "00000", "00000", "01111", "01111", "00001", "00001", "00001",
        "00001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "00001",
        "00001", "01111", "01111", "00001", "01111", "01111", "01111", "01111", "00001", "01111", "01111", "00001",
        "00001", "01111", "01111", "00001", "01111", "01111", "01111", "01111", "00001", "01111", "01111", "00001",
        "00001", "01111", "00001", "00001", "01111", "00001", "00001", "01111", "00001", "00001", "01111", "00001",
        "00001", "00001", "00001", "00001", "01111", "00001", "00001", "01111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "00001", "00001", "01111", "01111", "00001", "00001", "00001",
        -- 19
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "00001", "00001", "01111", "01111", "00001", "00001", "00001",
        "00001", "00001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "00001", "00001",
        "00001", "00001", "01111", "01111", "00110", "01111", "01111", "00110", "01111", "01111", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "01111", "01111", "01111", "01111", "00001", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "00110", "00110", "01111", "01111", "00001", "00001", "00001",
        "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111",
        "01111", "01111", "01111", "00001", "01111", "01111", "01111", "01111", "00001", "01111", "01111", "01111",
        "01111", "01111", "01111", "00001", "01111", "01111", "01111", "01111", "00001", "01111", "01111", "01111",
        "01111", "01111", "00001", "00001", "01111", "00001", "00001", "01111", "00001", "00001", "01111", "01111",
        "00001", "00001", "00001", "00001", "01111", "00001", "00001", "01111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "00001", "00001", "01111", "01111", "00001", "00001", "00001",
        -- 20
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "00001", "00001", "01111", "01111", "00001", "00001", "00001",
        "00001", "00001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "00001", "00001",
        "00001", "00001", "01111", "01111", "10010", "01111", "01111", "10010", "01111", "01111", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "01111", "01111", "01111", "01111", "00001", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "10010", "10010", "01111", "01111", "00001", "00001", "00001",
        "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111",
        "01111", "01111", "01111", "00001", "01111", "01111", "01111", "01111", "00001", "01111", "01111", "01111",
        "01111", "01111", "01111", "00001", "01111", "01111", "01111", "01111", "00001", "01111", "01111", "01111",
        "01111", "01111", "00001", "00001", "01111", "00001", "00001", "01111", "00001", "00001", "01111", "01111",
        "00001", "00001", "00001", "00001", "01111", "00001", "00001", "01111", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "01111", "01111", "00001", "00001", "01111", "01111", "00001", "00001", "00001",
        -- 21
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00000", "00000", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00001", "00101", "00101", "00101", "00101", "00001", "00101", "00001", "00001",
        "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        -- 22
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00000", "00000", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00001", "00101", "00101", "00101", "00101", "00001", "00101", "00001", "00001",
        "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00001",
        -- 23
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00000", "00000", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00001", "00101", "00101", "00101", "00101", "00001", "00101", "00001", "00001",
        "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        -- 24
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00000", "00000", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001",
        "00001", "00001", "00101", "00001", "00101", "00101", "00101", "00101", "00001", "00101", "00001", "00001",
        "00001", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        -- 25
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 26
        "00001", "00001", "00001", "00001", "00001", "00001", "01000", "01000", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "01000", "01000", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00000", "00001", "00001", "00001", "00001", "00001",
        "00001", "00000", "00000", "00000", "00001", "00000", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        -- 27
        "00001", "00001", "00001", "00001", "00001", "00001", "01000", "01000", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "01000", "01000", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00001", "00001", "00001", "00001", "00001",
        "00001", "00000", "00001", "00001", "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00000", "00000", "01100", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        -- 28
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "01000", "01000", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "00001", "00001", "00001",
        "00001", "00001", "00001", "00000", "00000", "00001", "01000", "01000", "00001", "00001", "00001", "00001",
        "00001", "00001", "00000", "00001", "00001", "00000", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        -- 29
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "01000", "01000", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "01000", "01000", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01000", "01000", "01000", "01000", "00001", "00001", "00001",
        "00001", "00001", "00000", "00001", "00001", "00001", "01000", "01000", "00001", "00001", "00001", "00001",
        "00001", "00000", "00001", "00000", "00001", "00000", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        -- 30
        "00001", "00001", "00001", "00001", "00001", "00001", "01010", "01010", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "01010", "01010", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00000", "00001", "00001", "00001", "00001", "00001",
        "00001", "00000", "00000", "00000", "00001", "00000", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        -- 31
        "00001", "00001", "00001", "00001", "00001", "00001", "01010", "01010", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "01010", "01010", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00001", "00001", "00001", "00001", "00001",
        "00001", "00000", "00001", "00001", "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00000", "00000", "01100", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        -- 32
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "01010", "01010", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "00001", "00001", "00001",
        "00001", "00001", "00001", "00000", "00000", "00001", "01010", "01010", "00001", "00001", "00001", "00001",
        "00001", "00001", "00000", "00001", "00001", "00000", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        -- 33
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "01010", "01010", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "01010", "01010", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "01010", "01010", "01010", "01010", "00001", "00001", "00001",
        "00001", "00001", "00000", "00001", "00001", "00001", "01010", "01010", "00001", "00001", "00001", "00001",
        "00001", "00000", "00001", "00000", "00001", "00000", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        -- 34
        "00011", "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00000", "00011", "00011", "00011", "00011", "00011",
        "00011", "00000", "00000", "00000", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00000", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 35
        "00011", "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00000", "00000", "00011", "00011", "00011", "00011", "00011",
        "00011", "00000", "00011", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00000", "00000", "01100", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 36
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00000", "00000", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00000", "00011", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 37
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00000", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00000", "00011", "00000", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00000", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 38
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 39
        "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010",
        "01010", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "01010",
        "01010", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "01010",
        "01010", "00001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "00001", "01010",
        "01010", "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001", "01010",
        "01010", "00001", "00001", "00101", "00101", "00000", "00000", "00101", "00101", "00001", "00001", "01010",
        "01010", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "01010",
        "01010", "00001", "00101", "00001", "00101", "00101", "00101", "00101", "00001", "00101", "00001", "01010",
        "01010", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "01010",
        "01010", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "01010",
        "01010", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "01010",
        "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010",
        -- 40
        "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010",
        "01010", "00001", "00001", "00111", "00111", "00001", "00001", "00111", "00111", "00001", "00001", "01010",
        "01010", "00001", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "00001", "01010",
        "01010", "00001", "00111", "00111", "00000", "00111", "00111", "00000", "00111", "00111", "00001", "01010",
        "01010", "00001", "00001", "00111", "00111", "00111", "00111", "00111", "00111", "00001", "01000", "01010",
        "01010", "00001", "00001", "00111", "00111", "00000", "00000", "00111", "00111", "00001", "00001", "01010",
        "01010", "00001", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00001", "01010",
        "01010", "00001", "00111", "00001", "00111", "00111", "00111", "00111", "00001", "00111", "00001", "01010",
        "01010", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00001", "00001", "00001", "01010",
        "01010", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00001", "00001", "00001", "01010",
        "01010", "00001", "00001", "00001", "00111", "00001", "00001", "00111", "00001", "00001", "00001", "01010",
        "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010",
        -- 41
        "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010",
        "01010", "00001", "01011", "00110", "00110", "01110", "01011", "00110", "00110", "01110", "00001", "01010",
        "01010", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "01010",
        "01010", "01011", "00110", "00110", "00000", "00110", "00110", "00000", "00110", "00110", "01110", "01010",
        "01010", "00001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "00001", "01010",
        "01010", "00001", "01011", "00110", "00110", "00000", "00000", "00110", "00110", "01110", "00001", "01010",
        "01010", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "01010",
        "01010", "01011", "00110", "01011", "00110", "00110", "00110", "00110", "01110", "00110", "01110", "01010",
        "01010", "00001", "01110", "00001", "00110", "00001", "00001", "00110", "00001", "01011", "00001", "01010",
        "01010", "00001", "00001", "00001", "00110", "00001", "00001", "00110", "00001", "00001", "00001", "01010",
        "01010", "00001", "00001", "00001", "01101", "00001", "00001", "01101", "00001", "00001", "00001", "01010",
        "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010",
        -- 42
        "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010",
        "01010", "00001", "00001", "10000", "10001", "00001", "00001", "10001", "10000", "00001", "00001", "01010",
        "01010", "00001", "10000", "00100", "10001", "10001", "10001", "10001", "00100", "10000", "00001", "01010",
        "01010", "00001", "10001", "10001", "00000", "10001", "10001", "00000", "10001", "10001", "00001", "01010",
        "01010", "00001", "00001", "10001", "10001", "10001", "10001", "10001", "10001", "00001", "00001", "01010",
        "01010", "00001", "00001", "10001", "10001", "00000", "00000", "10001", "10001", "00001", "00001", "01010",
        "01010", "00001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "00001", "01010",
        "01010", "00001", "10001", "00001", "10001", "10001", "10001", "10001", "00001", "10001", "00001", "01010",
        "01010", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "01010",
        "01010", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "01010",
        "01010", "00001", "00001", "00001", "10001", "00001", "00001", "10001", "00001", "00001", "00001", "01010",
        "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010",
        -- 43
        "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010",
        "01010", "00001", "00001", "01111", "01111", "00001", "00001", "01111", "01111", "00001", "00001", "01010",
        "01010", "00001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "00001", "01010",
        "01010", "00001", "01111", "01111", "00000", "01111", "01111", "00000", "01111", "01111", "00001", "01010",
        "01010", "00001", "00001", "01111", "01111", "01111", "01111", "01111", "01111", "00001", "00001", "01010",
        "01010", "00001", "00001", "01111", "01111", "00000", "00000", "01111", "01111", "00001", "00001", "01010",
        "01010", "00001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "00001", "01010",
        "01010", "00001", "01111", "00001", "01111", "01111", "01111", "01111", "00001", "01111", "00001", "01010",
        "01010", "00001", "00001", "00001", "01111", "00001", "00001", "01111", "00001", "00001", "00001", "01010",
        "01010", "00001", "00001", "00001", "01111", "00001", "00001", "01111", "00001", "00001", "00001", "01010",
        "01010", "00001", "00001", "00001", "01111", "00001", "00001", "01111", "00001", "00001", "00001", "01010",
        "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010",
        -- 44
        "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010",
        "01010", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "01010",
        "01010", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "01010",
        "01010", "00001", "00001", "00101", "00101", "00001", "00001", "00101", "00101", "00001", "00001", "01010",
        "01010", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "01010",
        "01010", "00001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "00001", "01010",
        "01010", "00001", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "00001", "01010",
        "01010", "00001", "00001", "00101", "00101", "00000", "00000", "00101", "00101", "00001", "00001", "01010",
        "01010", "00001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00001", "01010",
        "01010", "00001", "00101", "00001", "00101", "00101", "00101", "00101", "00001", "00101", "00001", "01010",
        "01010", "00001", "00001", "00001", "00101", "00001", "00001", "00101", "00001", "00001", "00001", "01010",
        "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010", "01010",
        -- 45
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
        "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
        "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
        "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00000", "00000",
        "00000", "00000", "00100", "00100", "00100", "00100", "00000", "00000", "00000", "00100", "00100", "00100",
        "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
        "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00000", "00000",
        "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
        "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
        "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 46
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100",
        "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100",
        "00100", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000", "00000", "00100", "00100",
        "00000", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00000",
        "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100",
        "00100", "00000", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00100",
        "00000", "00000", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00000",
        "00100", "00000", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00100",
        "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100",
        "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 47
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00100", "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00100", "00000", "00000",
        "00100", "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00100", "00000", "00000",
        "00100", "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00100", "00000", "00000",
        "00000", "00000", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00100", "00000", "00000",
        "00100", "00100", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000",
        "00100", "00100", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000",
        "00100", "00100", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000",
        "00100", "00100", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000",
        "00100", "00100", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 48
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "10010", "10010", "10010", "10010", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000",
        "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000",
        "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000",
        "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000",
        "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000",
        "00000", "00000", "10010", "00000", "00000", "00000", "10010", "00000", "00000", "10010", "00000", "00000",
        "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "10010", "00000", "00000",
        "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "10010", "10010", "10010", "10010", "00000", "10010", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 49
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "10010", "10010", "10010",
        "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
        "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
        "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
        "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
        "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
        "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
        "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
        "00000", "10010", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000", "10010",
        "00000", "00000", "10010", "10010", "10010", "00000", "00000", "00000", "00000", "10010", "10010", "10010",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 50
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "10010", "10010", "00000", "00000", "10010", "10010", "10010", "10010", "10010", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
        "10010", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 51
        "01110", "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110", "01110",
        "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110",
        "01110", "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110", "01110"
    );

    SIGNAL palette_index : unsigned(4 DOWNTO 0); -- max 32 colors
    SIGNAL full_color : STD_LOGIC_VECTOR(23 DOWNTO 0);
BEGIN
    -- get palette index from memory
    PROCESS (clk) BEGIN
        IF rising_edge(clk) THEN
            palette_index <= tile_rom_data(to_integer(address));
        END IF;
    END PROCESS;

    PROCESS (clk) BEGIN
        IF rising_edge(clk) THEN
            full_color <= palette_rom(to_integer(palette_index));
        END IF;
    END PROCESS;

    -- grab the high 4 bits of each color channel
    data_out <= full_color(23 DOWNTO 20) & full_color(15 DOWNTO 12) & full_color(7 DOWNTO 4);

END ARCHITECTURE;