LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY pMem IS
    PORT (
        adress : IN unsigned(11 DOWNTO 0);
        data : OUT STD_LOGIC_VECTOR(23 DOWNTO 0));
END pMem;

ARCHITECTURE func OF pMem IS
    TYPE p_mem_t IS ARRAY(NATURAL RANGE <>) OF STD_LOGIC_VECTOR(23 DOWNTO 0);
    CONSTANT p_mem_c : p_mem_t :=
    -- 00000_000_00_00_000000000000
    -- OP    GRx M  *  ADR 
    -- 5     3   2  2  12  
    (
    b"00000_101_00_00_000000000011", -- LOAD GR0, immediate, 0d60
    b"00000_000_00_00_000000000000", -- STORE 0
    b"00000_000_00_00_000000000010",
    b"00000_000_00_00_000000000100",
    b"00000_000_00_00_000000001000",
    b"00000_000_00_00_000000010000",
    b"00000_000_00_00_000000100000",
    b"00000_000_00_00_000010000000",
    b"00000_000_00_00_000000000000"
    );
BEGIN
    data <= p_mem_c(TO_INTEGER(adress));
END ARCHITECTURE;