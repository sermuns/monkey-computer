LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

-- usage: 
-- give uAddr, get uData at that address
ENTITY uMem IS
    PORT (
        address : IN unsigned(7 DOWNTO 0);
        data : OUT STD_LOGIC_VECTOR(22 DOWNTO 0));
END uMem;

ARCHITECTURE func OF uMem IS
    TYPE u_mem_t IS ARRAY(NATURAL RANGE <>) OF STD_LOGIC_VECTOR(22 DOWNTO 0);
    CONSTANT u_mem_array : u_mem_t :=
    -- 000_000_0000_0_0000_00000000
    -- TB _FB _ALU _P_SEQ _uADR
    (
    -- H�MTFAS
    b"010_000_0000_0_0000_00000000", --ASR := PC
    b"001_100_0000_1_0000_00000000", --IR := PM, PC++
    b"000_000_0000_0_0010_00000000", --uPC := K2

    -- ADDRESSERINGSFAS
    b"100_000_0000_0_0001_00000000", --ASR := IR, uPC := K1 (direkt)

    b"010_000_0000_1_0001_00000000", --ASR := PC, PC++, uPC:= K1 (omedelbar)
    b"100_000_0000_0_0000_00000000", --ASR := IR

    b"001_000_0000_0_0001_00000000", --ASR:= PM, uPC:= K1 (indirekt)

    b"100_011_0100_0_0000_00000000", --AR := IR (indexerad)
    b"101_011_0001_0_0000_00000000", --AR += GR3 (GR3 styrs av M)
    b"011_000_0000_0_0001_00000000", --ASR := AR, uPC := K1

    -- EXEKVERINGSFAS
    b"000_000_0000_0_0000_00000000",
    b"000_000_0000_0_0000_00000000",
    b"000_000_0000_0_0000_00000000",
    b"000_000_0000_0_0000_00000000",
    b"000_000_0000_0_0000_00000000",
    b"000_000_0000_0_0000_00000000",
    b"000_000_0000_0_0000_00000000",
    b"000_000_0000_0_0000_00000000",
    b"000_000_0000_0_0000_00000000",
    b"000_000_0000_0_0000_00000000",
    b"000_000_0000_0_0000_00000000",
    b"000_000_0000_0_0000_00000000"
    );
BEGIN
    data <= u_mem_array(TO_INTEGER(address));
END ARCHITECTURE;