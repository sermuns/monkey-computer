LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY pMem IS
    PORT (
        pAddr : IN unsigned(11 DOWNTO 0);
        pData : OUT unsigned(23 DOWNTO 0));
END pMem;

ARCHITECTURE func OF pMem IS
    TYPE p_mem_t IS ARRAY(11 DOWNTO 0) OF unsigned(23 DOWNTO 0);
    CONSTANT p_mem_c : p_mem_t :=
    --"00000_000_00_00000000000000" = "OP_GRx_M_ADR"
    (
    b"00001_000_00_00000000000000",
    b"00000_000_00_10000000000000",
    b"00000_000_00_00000000000000",
    b"00000_000_00_10000000000000",
    b"00000_000_00_10000000000000",
    b"00000_000_00_10000000000000",
    b"00000_000_00_10000000000000",
    b"00000_000_00_00000000000000",
    b"00000_000_00_00000000000000",
    b"00000_000_00_00000000000000",
    b"00000_000_00_00000000000000",
    b"00000_000_00_00000000000000",
    b"00000_000_00_00000000000000",
    b"00000_000_00_00000000000000",
    b"00000_000_00_00000000000000",
    b"00000_000_00_00000000000000"
    );

    SIGNAL p_mem : p_mem_t := p_mem_c;

BEGIN
    pData <= p_mem(TO_INTEGER(pAddr));
END ARCHITECTURE;