LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY tile_rom IS
    PORT (
        clk : IN STD_LOGIC;
        address : IN UNSIGNED(13 DOWNTO 0); -- 14 bit address
        data_out : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
    );
END tile_rom;

ARCHITECTURE func OF tile_rom IS TYPE palette_rom_type IS ARRAY(0 TO 18) OF STD_LOGIC_VECTOR(23 DOWNTO 0);
    CONSTANT palette_rom : palette_rom_type := (
        00 => x"000000",
        01 => x"ffffff",
        02 => x"332222",
        03 => x"404040",
        04 => x"f5a097",
        05 => x"774433",
        06 => x"993311",
        07 => x"cc8855",
        08 => x"ffdd55",
        09 => x"176b04",
        10 => x"44eebb",
        11 => x"3388dd",
        12 => x"070708",
        13 => x"555577",
        14 => x"5544aa",
        15 => x"422433",
        16 => x"73172d",
        17 => x"e86a73",
        18 => x"b4202a"
    );
    CONSTANT TILE_SIZE : INTEGER := 12 * 12;

    TYPE tile_rom_type IS ARRAY(0 TO 9359) OF unsigned(4 DOWNTO 0);
    CONSTANT tile_rom_data : tile_rom_type := (
        -- 0
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        -- 1
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00000", "00000", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "01001", "00101", "00101", "00101", "00101", "01001", "00101", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        -- 2
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00000", "00000", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "01001", "00101", "00101", "00101", "00101", "01001", "00101", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        -- 3
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00000", "00000", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "01001", "00101", "00101", "00101", "00101", "01001", "00101", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        -- 4
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00000", "00000", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "01001", "00101", "00101", "00101", "00101", "01001", "00101", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        -- 5
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00111", "00111", "01001", "01001", "00111", "00111", "01001", "01001", "01001",
        "01001", "01001", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "01001", "01001",
        "01001", "01001", "00111", "00111", "00000", "00111", "00111", "00000", "00111", "00111", "01001", "01001",
        "01001", "01001", "01001", "00111", "00111", "00111", "00111", "00111", "00111", "01001", "01000", "01001",
        "01001", "01001", "01001", "00111", "00111", "00000", "00000", "00111", "00111", "01001", "01001", "01001",
        "01001", "01001", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "01001", "01001",
        "01001", "01001", "00111", "01001", "00111", "00111", "00111", "00111", "01001", "00111", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00111", "00111", "01001", "01001", "00111", "00111", "01001", "01001", "01001",
        -- 6
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00111", "00111", "01001", "01001", "00111", "00111", "01001", "01001", "01001",
        "01001", "01001", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "01001", "01001",
        "01001", "01001", "00111", "00111", "00000", "00111", "00111", "00000", "00111", "00111", "01001", "01001",
        "01001", "01001", "01001", "00111", "00111", "00111", "00111", "00111", "00111", "01001", "01000", "01001",
        "01001", "01001", "01001", "00111", "00111", "00000", "00000", "00111", "00111", "01001", "01001", "01001",
        "01001", "01001", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "01001", "01001",
        "01001", "01001", "00111", "01001", "00111", "00111", "00111", "00111", "01001", "00111", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "00111", "01001", "01001", "01001",
        "01001", "01001", "01001", "00111", "00111", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        -- 7
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00111", "00111", "01001", "01001", "00111", "00111", "01001", "01001", "01001",
        "01001", "01001", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "01001", "01001",
        "01001", "01001", "00111", "00111", "00000", "00111", "00111", "00000", "00111", "00111", "01001", "01001",
        "01001", "01001", "01001", "00111", "00111", "00111", "00111", "00111", "00111", "01001", "01000", "01001",
        "01001", "01001", "01001", "00111", "00111", "00000", "00000", "00111", "00111", "01001", "01001", "01001",
        "01001", "01001", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "01001", "01001",
        "01001", "01001", "00111", "01001", "00111", "00111", "00111", "00111", "01001", "00111", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00111", "00111", "01001", "01001", "00111", "00111", "01001", "01001", "01001",
        -- 8
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00111", "00111", "01001", "01001", "00111", "00111", "01001", "01001", "01001",
        "01001", "01001", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "01001", "01001",
        "01001", "01001", "00111", "00111", "00000", "00111", "00111", "00000", "00111", "00111", "01001", "01001",
        "01001", "01001", "01001", "00111", "00111", "00111", "00111", "00111", "00111", "01001", "01000", "01001",
        "01001", "01001", "01001", "00111", "00111", "00000", "00000", "00111", "00111", "01001", "01001", "01001",
        "01001", "01001", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "01001", "01001",
        "01001", "01001", "00111", "01001", "00111", "00111", "00111", "00111", "01001", "00111", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "00111", "01001", "01001", "01001",
        "01001", "01001", "01001", "00111", "00111", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        -- 9
        "01001", "01001", "01001", "01110", "01011", "01001", "01001", "01110", "01011", "01001", "01001", "01001",
        "01001", "01001", "01011", "00110", "00110", "01110", "01011", "00110", "00110", "01110", "01001", "01001",
        "01001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "01001",
        "01001", "01011", "00110", "00110", "00000", "00110", "00110", "00000", "00110", "00110", "01110", "01001",
        "01001", "01001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "01001", "01001",
        "01001", "01001", "01011", "00110", "00110", "00000", "00000", "00110", "00110", "01110", "01001", "01001",
        "01001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "01001",
        "01001", "01011", "00110", "01011", "00110", "00110", "00110", "00110", "01110", "00110", "01110", "01001",
        "01001", "01001", "01110", "01001", "00110", "01001", "01001", "00110", "01001", "01011", "01001", "01001",
        "01001", "01001", "01001", "01001", "00110", "01001", "01001", "00110", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01101", "01001", "01001", "01101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01101", "01101", "01001", "01001", "01101", "01101", "01001", "01001", "01001",
        -- 10
        "01001", "01001", "01001", "01011", "01110", "01001", "01001", "01011", "01110", "01001", "01001", "01001",
        "01001", "01001", "01110", "00110", "00110", "01011", "01110", "00110", "00110", "01011", "01001", "01001",
        "01001", "01011", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01110", "01001",
        "01001", "01110", "00110", "00110", "00000", "00110", "00110", "00000", "00110", "00110", "01011", "01001",
        "01001", "01001", "01011", "00110", "00110", "00110", "00110", "00110", "00110", "01110", "01001", "01001",
        "01001", "01001", "01110", "00110", "00110", "00000", "00000", "00110", "00110", "01011", "01001", "01001",
        "01001", "01011", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01110", "01001",
        "01001", "01110", "00110", "01110", "00110", "00110", "00110", "00110", "01011", "00110", "01011", "01001",
        "01001", "01001", "01011", "01001", "00110", "01001", "01001", "00110", "01001", "01110", "01001", "01001",
        "01001", "01001", "01001", "01001", "00110", "01001", "01001", "00110", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01101", "01001", "01001", "01101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01101", "01101", "01001", "01001", "01101", "01101", "01001", "01001", "01001",
        -- 11
        "01001", "01001", "01001", "01110", "01011", "01001", "01001", "01110", "01011", "01001", "01001", "01001",
        "01001", "01001", "01011", "00110", "00110", "01110", "01011", "00110", "00110", "01110", "01001", "01001",
        "01001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "01001",
        "01001", "01011", "00110", "00110", "00000", "00110", "00110", "00000", "00110", "00110", "01110", "01001",
        "01001", "01001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "01001", "01001",
        "01001", "01001", "01011", "00110", "00110", "00000", "00000", "00110", "00110", "01110", "01001", "01001",
        "01001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "01001",
        "01001", "01011", "00110", "01011", "00110", "00110", "00110", "00110", "01110", "00110", "01110", "01001",
        "01001", "01001", "01110", "01001", "00110", "01001", "01001", "00110", "01001", "01011", "01001", "01001",
        "01001", "01001", "01001", "01001", "00110", "01001", "01001", "00110", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01101", "01001", "01001", "01101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01101", "01101", "01001", "01001", "01101", "01101", "01001", "01001", "01001",
        -- 12
        "01001", "01001", "01001", "01011", "01110", "01001", "01001", "01011", "01110", "01001", "01001", "01001",
        "01001", "01001", "01110", "00110", "00110", "01011", "01110", "00110", "00110", "01011", "01001", "01001",
        "01001", "01011", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01110", "01001",
        "01001", "01110", "00110", "00110", "00000", "00110", "00110", "00000", "00110", "00110", "01011", "01001",
        "01001", "01001", "01011", "00110", "00110", "00110", "00110", "00110", "00110", "01110", "01001", "01001",
        "01001", "01001", "01110", "00110", "00110", "00000", "00000", "00110", "00110", "01011", "01001", "01001",
        "01001", "01011", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01110", "01001",
        "01001", "01110", "00110", "01110", "00110", "00110", "00110", "00110", "01011", "00110", "01011", "01001",
        "01001", "01001", "01011", "01001", "00110", "01001", "01001", "00110", "01001", "01110", "01001", "01001",
        "01001", "01001", "01001", "01001", "00110", "01001", "01001", "00110", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01101", "01001", "01001", "01101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01101", "01101", "01001", "01001", "01101", "01101", "01001", "01001", "01001",
        -- 13
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "10000", "10001", "01001", "01001", "10001", "10000", "01001", "01001", "01001",
        "01001", "01001", "10000", "00100", "10001", "10001", "10001", "10001", "00100", "10000", "01001", "01001",
        "01001", "01001", "10001", "10001", "00000", "10001", "10001", "00000", "10001", "10001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "10001", "10001", "10001", "10001", "01001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "00000", "00000", "10001", "10001", "01001", "01001", "01001",
        "01001", "01001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "01001", "01001",
        "01001", "01001", "10001", "01001", "10001", "10001", "10001", "10001", "01001", "10001", "01001", "01001",
        "01001", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "01001", "01001", "10001", "10001", "01001", "01001", "01001",
        -- 14
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "10000", "10001", "01001", "01001", "10001", "10000", "01001", "01001", "01001",
        "01001", "01001", "10000", "00100", "10001", "10001", "10001", "10001", "00100", "10000", "01001", "01001",
        "01001", "01001", "10001", "10001", "00000", "10001", "10001", "00000", "10001", "10001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "10001", "10001", "10001", "10001", "01001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "00000", "00000", "10001", "10001", "01001", "01001", "01001",
        "01001", "01001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "01001", "01001",
        "01001", "01001", "10001", "01001", "10001", "10001", "10001", "10001", "01001", "10001", "01001", "01001",
        "01001", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "10001", "01001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        -- 15
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "10000", "10001", "01001", "01001", "10001", "10000", "01001", "01001", "01001",
        "01001", "01001", "10000", "00100", "10001", "10001", "10001", "10001", "00100", "10000", "01001", "01001",
        "01001", "01001", "10001", "10001", "00000", "10001", "10001", "00000", "10001", "10001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "10001", "10001", "10001", "10001", "01001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "00000", "00000", "10001", "10001", "01001", "01001", "01001",
        "01001", "01001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "01001", "01001",
        "01001", "01001", "10001", "01001", "10001", "10001", "10001", "10001", "01001", "10001", "01001", "01001",
        "01001", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "01001", "01001", "10001", "10001", "01001", "01001", "01001",
        -- 16
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "10000", "10001", "01001", "01001", "10001", "10000", "01001", "01001", "01001",
        "01001", "01001", "10000", "00100", "10001", "10001", "10001", "10001", "00100", "10000", "01001", "01001",
        "01001", "01001", "10001", "10001", "00000", "10001", "10001", "00000", "10001", "10001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "10001", "10001", "10001", "10001", "01001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "00000", "00000", "10001", "10001", "01001", "01001", "01001",
        "01001", "01001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "01001", "01001",
        "01001", "01001", "10001", "01001", "10001", "10001", "10001", "10001", "01001", "10001", "01001", "01001",
        "01001", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "10001", "10001", "01001", "01001", "01001",
        -- 17
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "01001", "01001", "01111", "01111", "01001", "01001", "01001",
        "01001", "01001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01001", "01001",
        "01001", "01001", "01111", "01111", "00000", "01111", "01111", "00000", "01111", "01111", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "01111", "01111", "01111", "01111", "01001", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "00000", "00000", "01111", "01111", "01001", "01001", "01001",
        "01001", "01001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01001", "01001",
        "01001", "01001", "01111", "01001", "01111", "01111", "01111", "01111", "01001", "01111", "01001", "01001",
        "01001", "01001", "01001", "01001", "01111", "01001", "01001", "01111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01111", "01001", "01001", "01111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01111", "01001", "01001", "01111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "01001", "01001", "01111", "01111", "01001", "01001", "01001",
        -- 18
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "01001", "01001", "01111", "01111", "01001", "01001", "01001",
        "01001", "01001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01001", "01001",
        "01001", "01001", "01111", "01111", "00000", "01111", "01111", "00000", "01111", "01111", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "01111", "01111", "01111", "01111", "01001", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "00000", "00000", "01111", "01111", "01001", "01001", "01001",
        "01001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01001",
        "01001", "01111", "01111", "01001", "01111", "01111", "01111", "01111", "01001", "01111", "01111", "01001",
        "01001", "01111", "01111", "01001", "01111", "01111", "01111", "01111", "01001", "01111", "01111", "01001",
        "01001", "01111", "01001", "01001", "01111", "01001", "01001", "01111", "01001", "01001", "01111", "01001",
        "01001", "01001", "01001", "01001", "01111", "01001", "01001", "01111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "01001", "01001", "01111", "01111", "01001", "01001", "01001",
        -- 19
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "01001", "01001", "01111", "01111", "01001", "01001", "01001",
        "01001", "01001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01001", "01001",
        "01001", "01001", "01111", "01111", "00110", "01111", "01111", "00110", "01111", "01111", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "01111", "01111", "01111", "01111", "01001", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "00110", "00110", "01111", "01111", "01001", "01001", "01001",
        "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111",
        "01111", "01111", "01111", "01001", "01111", "01111", "01111", "01111", "01001", "01111", "01111", "01111",
        "01111", "01111", "01111", "01001", "01111", "01111", "01111", "01111", "01001", "01111", "01111", "01111",
        "01111", "01111", "01001", "01001", "01111", "01001", "01001", "01111", "01001", "01001", "01111", "01111",
        "01001", "01001", "01001", "01001", "01111", "01001", "01001", "01111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "01001", "01001", "01111", "01111", "01001", "01001", "01001",
        -- 20
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "01001", "01001", "01111", "01111", "01001", "01001", "01001",
        "01001", "01001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01001", "01001",
        "01001", "01001", "01111", "01111", "10010", "01111", "01111", "10010", "01111", "01111", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "01111", "01111", "01111", "01111", "01001", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "10010", "10010", "01111", "01111", "01001", "01001", "01001",
        "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111",
        "01111", "01111", "01111", "01001", "01111", "01111", "01111", "01111", "01001", "01111", "01111", "01111",
        "01111", "01111", "01111", "01001", "01111", "01111", "01111", "01111", "01001", "01111", "01111", "01111",
        "01111", "01111", "01001", "01001", "01111", "01001", "01001", "01111", "01001", "01001", "01111", "01111",
        "01001", "01001", "01001", "01001", "01111", "01001", "01001", "01111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "01001", "01001", "01111", "01111", "01001", "01001", "01001",
        -- 21
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00000", "00000", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "01001", "00101", "00101", "00101", "00101", "01001", "00101", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        -- 22
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00000", "00000", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "01001", "00101", "00101", "00101", "00101", "01001", "00101", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "01001", "01001", "01001", "01001", "00101", "01001", "01001", "01001",
        -- 23
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00000", "00000", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "01001", "00101", "00101", "00101", "00101", "01001", "00101", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        -- 24
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00000", "00000", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "01001", "00101", "00101", "00101", "00101", "01001", "00101", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        -- 25
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 26
        "00011", "00011", "00011", "00011", "00011", "00011", "01000", "01000", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "01000", "01000", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00000", "00011", "00011", "00011", "00011", "00011",
        "00011", "00000", "00000", "00000", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00000", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 27
        "00011", "00011", "00011", "00011", "00011", "00011", "01000", "01000", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "01000", "01000", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00000", "00000", "00011", "00011", "00011", "00011", "00011",
        "00011", "00000", "00011", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00000", "00000", "01100", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 28
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "01000", "01000", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "00011", "00011", "00011",
        "00011", "00011", "00011", "00000", "00000", "00011", "01000", "01000", "00011", "00011", "00011", "00011",
        "00011", "00011", "00000", "00011", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 29
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "01000", "01000", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "01000", "01000", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01000", "01000", "01000", "01000", "00011", "00011", "00011",
        "00011", "00011", "00000", "00011", "00011", "00011", "01000", "01000", "00011", "00011", "00011", "00011",
        "00011", "00000", "00011", "00000", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00000", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 30
        "00011", "00011", "00011", "00011", "00011", "00011", "01010", "01010", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "01010", "01010", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00000", "01001", "00011", "00011", "00011", "00011",
        "00011", "00000", "00000", "00000", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00000", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 31
        "00011", "00011", "00011", "00011", "00011", "00011", "01010", "01010", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "01010", "01010", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00000", "00000", "00011", "00011", "00011", "00011", "00011",
        "00011", "00000", "00011", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00000", "00000", "01100", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 32
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "01010", "01010", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "00011", "00011", "00011",
        "00011", "00011", "00011", "00000", "00000", "00011", "01010", "01010", "00011", "00011", "00011", "00011",
        "00011", "00011", "00000", "00011", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 33
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "01010", "01010", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "01010", "01010", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "01010", "01010", "01010", "01010", "00011", "00011", "00011",
        "00011", "00011", "00000", "00011", "00011", "00011", "01010", "01010", "00011", "00011", "00011", "00011",
        "00011", "00000", "00011", "00000", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00000", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 34
        "00011", "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00000", "00011", "00011", "00011", "00011", "00011",
        "00011", "00000", "00000", "00000", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00000", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 35
        "00011", "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00000", "00000", "00011", "00011", "00011", "00011", "00011",
        "00011", "00000", "00011", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00000", "00000", "01100", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 36
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00000", "00000", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00000", "00011", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 37
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00111", "00111", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00111", "00111", "00111", "00111", "00011", "00011", "00011",
        "00011", "00011", "00000", "00011", "00011", "00011", "00111", "00111", "00011", "00011", "00011", "00011",
        "00011", "00000", "00011", "00000", "00011", "00000", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00000", "00000", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        -- 38
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 39
        "01110", "01110", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01110", "01110",
        "01110", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01110",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00000", "00000", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "01001", "00101", "00101", "00101", "00101", "01001", "00101", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01001",
        "01110", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01110",
        "01110", "01110", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01110", "01110",
        -- 40
        "01110", "01110", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01110", "01110",
        "01110", "01001", "01001", "00111", "00111", "01001", "01001", "00111", "00111", "01001", "01001", "01110",
        "01001", "01001", "00111", "00010", "00010", "00010", "00010", "00010", "00010", "00111", "01001", "01001",
        "01001", "01001", "00111", "00111", "00000", "00111", "00111", "00000", "00111", "00111", "01001", "01001",
        "01001", "01001", "01001", "00111", "00111", "00111", "00111", "00111", "00111", "01001", "01000", "01001",
        "01001", "01001", "01001", "00111", "00111", "00000", "00000", "00111", "00111", "01001", "01001", "01001",
        "01001", "01001", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "00111", "01001", "01001",
        "01001", "01001", "00111", "01001", "00111", "00111", "00111", "00111", "01001", "00111", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "01001", "01001", "01001", "01001",
        "01110", "01001", "01001", "01001", "00111", "01001", "01001", "00111", "01001", "01001", "01001", "01110",
        "01110", "01110", "01001", "00111", "00111", "01001", "01001", "00111", "00111", "01001", "01110", "01110",
        -- 41
        "01110", "01110", "01001", "01110", "01011", "01001", "01001", "01110", "01011", "01001", "01110", "01110",
        "01110", "01001", "01011", "00110", "00110", "01110", "01011", "00110", "00110", "01110", "01001", "01110",
        "01001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "01001",
        "01001", "01011", "00110", "00110", "00000", "00110", "00110", "00000", "00110", "00110", "01110", "01001",
        "01001", "01001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "01001", "01001",
        "01001", "01001", "01011", "00110", "00110", "00000", "00000", "00110", "00110", "01110", "01001", "01001",
        "01001", "01110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "00110", "01011", "01001",
        "01001", "01011", "00110", "01011", "00110", "00110", "00110", "00110", "01110", "00110", "01110", "01001",
        "01001", "01001", "01110", "01001", "00110", "01001", "01001", "00110", "01001", "01011", "01001", "01001",
        "01001", "01001", "01001", "01001", "00110", "01001", "01001", "00110", "01001", "01001", "01001", "01001",
        "01110", "01001", "01001", "01001", "01101", "01001", "01001", "01101", "01001", "01001", "01001", "01110",
        "01110", "01110", "01001", "01101", "01101", "01001", "01001", "01101", "01101", "01001", "01110", "01110",
        -- 42
        "01110", "01110", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01110", "01110",
        "01110", "01001", "01001", "10000", "10001", "01001", "01001", "10001", "10000", "01001", "01001", "01110",
        "01001", "01001", "10000", "00100", "10001", "10001", "10001", "10001", "00100", "10000", "01001", "01001",
        "01001", "01001", "10001", "10001", "00000", "10001", "10001", "00000", "10001", "10001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "10001", "10001", "10001", "10001", "01001", "01001", "01001",
        "01001", "01001", "01001", "10001", "10001", "00000", "00000", "10001", "10001", "01001", "01001", "01001",
        "01001", "01001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "10001", "01001", "01001",
        "01001", "01001", "10001", "01001", "10001", "10001", "10001", "10001", "01001", "10001", "01001", "01001",
        "01001", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01001",
        "01110", "01001", "01001", "01001", "10001", "01001", "01001", "10001", "01001", "01001", "01001", "01110",
        "01110", "01110", "01001", "10001", "10001", "01001", "01001", "10001", "10001", "01001", "01110", "01110",
        -- 43
        "01110", "01110", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01110", "01110",
        "01110", "01001", "01001", "01111", "01111", "01001", "01001", "01111", "01111", "01001", "01001", "01110",
        "01001", "01001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01001", "01001",
        "01001", "01001", "01111", "01111", "00000", "01111", "01111", "00000", "01111", "01111", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "01111", "01111", "01111", "01111", "01001", "01001", "01001",
        "01001", "01001", "01001", "01111", "01111", "00000", "00000", "01111", "01111", "01001", "01001", "01001",
        "01001", "01001", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01111", "01001", "01001",
        "01001", "01001", "01111", "01001", "01111", "01111", "01111", "01111", "01001", "01111", "01001", "01001",
        "01001", "01001", "01001", "01001", "01111", "01001", "01001", "01111", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "01001", "01111", "01001", "01001", "01111", "01001", "01001", "01001", "01001",
        "01110", "01001", "01001", "01001", "01111", "01001", "01001", "01111", "01001", "01001", "01001", "01110",
        "01110", "01110", "01001", "01111", "01111", "01001", "01001", "01111", "01111", "01001", "01110", "01110",
        -- 44
        "01110", "01110", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01110", "01110",
        "01110", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01110",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "00101", "00000", "00101", "00101", "00000", "00101", "00101", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "01001", "00101", "00101", "00000", "00000", "00101", "00101", "01001", "01001", "01001",
        "01001", "01001", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "00101", "01001", "01001",
        "01001", "01001", "00101", "01001", "00101", "00101", "00101", "00101", "01001", "00101", "01001", "01001",
        "01110", "01001", "01001", "01001", "00101", "01001", "01001", "00101", "01001", "01001", "01001", "01110",
        "01110", "01110", "01001", "00101", "00101", "01001", "01001", "00101", "00101", "01001", "01110", "01110",
        -- 45
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00100", "00100", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00100", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 46
        "01110", "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110", "01110",
        "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110",
        "00000", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00100", "00100", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00100", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00000", "00000", "00000",
        "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00000", "00000", "00000",
        "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110",
        "01110", "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110", "01110",
        -- 47
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "10010", "10010", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "10010", "00000", "00000", "10010", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000",
        "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000",
        "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000",
        "00000", "00000", "00000", "10010", "00000", "00000", "10010", "00000", "10010", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "10010", "00000", "00000", "10010", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "10010", "10010", "00000", "10010", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 48
        "01110", "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110", "01110",
        "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110",
        "00000", "00000", "00000", "00000", "00000", "10010", "10010", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "10010", "00000", "00000", "10010", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000",
        "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000",
        "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000",
        "00000", "00000", "00000", "10010", "00000", "00000", "10010", "00000", "10010", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "10010", "00000", "00000", "10010", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "10010", "10010", "00000", "10010", "00000", "00000", "00000",
        "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110",
        "01110", "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110", "01110",
        -- 49
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "01010", "00000", "00000", "01010", "00000", "01010", "01010", "01010", "00000", "00000",
        "00000", "00000", "01010", "00000", "00000", "01010", "00000", "01010", "00000", "00000", "01010", "00000",
        "00000", "00000", "01010", "01010", "01010", "01010", "00000", "01010", "00000", "00000", "01010", "00000",
        "00000", "00000", "01010", "01010", "01010", "01010", "00000", "01010", "01010", "01010", "00000", "00000",
        "00000", "00000", "01010", "00000", "00000", "01010", "00000", "01010", "00000", "00000", "00000", "00000",
        "00000", "00000", "01010", "00000", "00000", "01010", "00000", "01010", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 50
        "01110", "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110", "01110",
        "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "01010", "00000", "00000", "01010", "00000", "01010", "01010", "01010", "00000", "00000",
        "00000", "00000", "01010", "00000", "00000", "01010", "00000", "01010", "00000", "00000", "01010", "00000",
        "00000", "00000", "01010", "01010", "01010", "01010", "00000", "01010", "00000", "00000", "01010", "00000",
        "00000", "00000", "01010", "01010", "01010", "01010", "00000", "01010", "01010", "01010", "00000", "00000",
        "00000", "00000", "01010", "00000", "00000", "01010", "00000", "01010", "00000", "00000", "00000", "00000",
        "00000", "00000", "01010", "00000", "00000", "01010", "00000", "01010", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110",
        "01110", "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110", "01110",
        -- 51
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "01000", "01000", "01000", "01000", "01000", "01000", "00000", "00000", "00000",
        "00000", "00000", "01000", "01000", "01000", "00000", "00000", "00000", "01000", "01000", "00000", "00000",
        "00000", "01000", "01000", "01000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "01000", "01000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "01000", "01000", "00000", "00000", "00000", "01000", "01000", "01000", "01000", "00000", "00000",
        "00000", "01000", "01000", "01000", "00000", "00000", "00000", "01000", "01000", "00000", "00000", "00000",
        "00000", "00000", "01000", "01000", "01000", "00000", "00000", "01000", "01000", "00000", "00000", "00000",
        "00000", "00000", "00000", "01000", "01000", "01000", "01000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 52
        "01110", "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110", "01110",
        "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110",
        "00000", "00000", "00000", "01000", "01000", "01000", "01000", "01000", "01000", "00000", "00000", "00000",
        "00000", "00000", "01000", "01000", "01000", "00000", "00000", "00000", "01000", "01000", "00000", "00000",
        "00000", "01000", "01000", "01000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "01000", "01000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "01000", "01000", "00000", "00000", "00000", "01000", "01000", "01000", "01000", "00000", "00000",
        "00000", "01000", "01000", "01000", "00000", "00000", "00000", "01000", "01000", "00000", "00000", "00000",
        "00000", "00000", "01000", "01000", "01000", "00000", "00000", "01000", "01000", "00000", "00000", "00000",
        "00000", "00000", "00000", "01000", "01000", "01000", "01000", "00000", "00000", "00000", "00000", "00000",
        "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110",
        "01110", "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110", "01110",
        -- 53
        "01110", "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110", "01110",
        "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110",
        "01110", "01110", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "01110", "01110",
        -- 54
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00001", "00000", "00000", "00001", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00001", "00000", "00000", "00001", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 55
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00001", "00001", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00001", "00001", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00001", "00001", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00001", "00001", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00001", "00001", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 56
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 57
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 58
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 59
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 60
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 61
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 62
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 63
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00001", "00000", "00000", "00000", "00000", "00001", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        -- 64
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000"
    );

    SIGNAL palette_index : unsigned(4 DOWNTO 0); -- max 32 colors
    SIGNAL full_color : STD_LOGIC_VECTOR(23 DOWNTO 0);
BEGIN
    -- get palette index from memory
    PROCESS (clk) BEGIN
        IF rising_edge(clk) THEN
            palette_index <= tile_rom_data(to_integer(address));
        END IF;
    END PROCESS;

    PROCESS (clk) BEGIN
        IF rising_edge(clk) THEN
            full_color <= palette_rom(to_integer(palette_index));
        END IF;
    END PROCESS;

    -- grab the high 4 bits of each color channel
    data_out <= full_color(23 DOWNTO 20) & full_color(15 DOWNTO 12) & full_color(7 DOWNTO 4);

END ARCHITECTURE;
