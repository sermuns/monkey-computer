LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY tile_rom_menu IS
    PORT (
        clk : IN STD_LOGIC;
        address : IN UNSIGNED(13 DOWNTO 0); -- 14 bit address
        menu_data_out : OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
    );
END tile_rom_menu;

ARCHITECTURE func_menu OF tile_rom_menu IS TYPE palette_rom_type IS ARRAY(0 TO 18) OF STD_LOGIC_VECTOR(23 DOWNTO 0);
    CONSTANT palette_rom : palette_rom_type := (
        00 => x"000000",
        01 => x"ffffff",
        02 => x"332222",
        03 => x"404040",
        04 => x"f5a097",
        05 => x"774433",
        06 => x"993311",
        07 => x"cc8855",
        08 => x"ffdd55",
        09 => x"176b04",
        10 => x"44eebb",
        11 => x"3388dd",
        12 => x"070708",
        13 => x"555577",
        14 => x"5544aa",
        15 => x"422433",
        16 => x"73172d",
        17 => x"e86a73",
        18 => x"b4202a"
    );
    CONSTANT TILE_SIZE : INTEGER := 12 * 12;

    TYPE tile_rom_menu_type IS ARRAY(0 TO 4000) OF unsigned(4 DOWNTO 0);
    CONSTANT tile_rom_menu_data : tile_rom_menu_type := (
        -- 0
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "01110", "01011", "00000", "00000", "01110", "01011", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00001", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "00000", "00000", "00000", "01110", "01011", "00000", "00000", "01110", "01011", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
        "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "01001", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
 
        -- RESET and QUIT ROM
                -- 45
                "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
                "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
                "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
                "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
                "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00000", "00000",
                "00000", "00000", "00100", "00100", "00100", "00100", "00000", "00000", "00000", "00100", "00100", "00100",
                "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
                "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00000", "00000",
                "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
                "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
                "00000", "00000", "00100", "00100", "00000", "00100", "00100", "00000", "00000", "00100", "00100", "00100",
                "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
                -- 46
                "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
                "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100",
                "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100",
                "00100", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000", "00000", "00100", "00100",
                "00000", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00000",
                "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100",
                "00100", "00000", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00100",
                "00000", "00000", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00000",
                "00100", "00000", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00100", "00100",
                "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100",
                "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00000", "00000", "00100", "00100",
                "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
                -- 47
                "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
                "00100", "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00100", "00000", "00000",
                "00100", "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00100", "00000", "00000",
                "00100", "00100", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00100", "00000", "00000",
                "00000", "00000", "00000", "00000", "00100", "00100", "00100", "00100", "00100", "00100", "00000", "00000",
                "00100", "00100", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000",
                "00100", "00100", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000",
                "00000", "00000", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000",
                "00100", "00100", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000",
                "00100", "00100", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000",
                "00100", "00100", "00000", "00000", "00000", "00000", "00100", "00100", "00000", "00000", "00000", "00000",
                "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
                -- 48
                "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
                "00000", "00000", "00000", "00000", "10010", "10010", "10010", "10010", "00000", "00000", "00000", "00000",
                "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000",
                "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000",
                "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000",
                "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000",
                "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000",
                "00000", "00000", "10010", "00000", "00000", "00000", "10010", "00000", "00000", "10010", "00000", "00000",
                "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "10010", "00000", "00000",
                "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000",
                "00000", "00000", "00000", "00000", "10010", "10010", "10010", "10010", "00000", "10010", "00000", "00000",
                "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
                -- 49
                "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
                "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "10010", "10010", "10010",
                "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
                "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
                "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
                "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
                "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
                "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
                "10010", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "10010",
                "00000", "10010", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000", "10010",
                "00000", "00000", "10010", "10010", "10010", "00000", "00000", "00000", "00000", "10010", "10010", "10010",
                "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
                -- 50
                "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",
                "10010", "10010", "00000", "00000", "10010", "10010", "10010", "10010", "10010", "00000", "00000", "00000",
                "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
                "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
                "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
                "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
                "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
                "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
                "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
                "00000", "00000", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
                "10010", "10010", "00000", "00000", "00000", "00000", "10010", "00000", "00000", "00000", "00000", "00000",
                "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000", "00000",

        OTHERS => (OTHERS => 'U')
    );

    SIGNAL palette_index : unsigned(4 DOWNTO 0); -- max 32 colors
BEGIN
    PROCESS (address)
    BEGIN
        -- get palette index from memory
        palette_index <= tile_rom_menu_data(to_integer(address));
        menu_data_out <= palette_rom(to_integer(palette_index));
    END PROCESS;
END ARCHITECTURE;