LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY tile_rom IS
    PORT (
        address : IN UNSIGNED(13 DOWNTO 0); -- 14 bit address
        data_out : OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
    );
END tile_rom;

ARCHITECTURE func OF tile_rom IS
    TYPE palette_rom_type IS ARRAY(0 TO 31) OF STD_LOGIC_VECTOR(23 DOWNTO 0);
    CONSTANT palette_rom : palette_rom_type := (
        0 => X"ffffff",
        1 => X"000000",
        2 => X"332222",
        3 => X"404040",
        4 => X"6c6c6c",
        5 => X"909090",
        6 => X"f5a097",
        7 => X"774433",
        8 => X"993311",
        9 => X"cc8855",
        10 => X"c89870",
        11 => X"dcac84",
        12 => X"b48458",
        13 => X"dd7711",
        14 => X"a08662",
        15 => X"ecd09c",
        16 => X"ffdd55",
        17 => X"2f6e1e",
        18 => X"1c6e09",
        19 => X"176b04",
        20 => X"114c04",
        21 => X"3eff30",
        22 => X"2bff44",
        23 => X"44eebb",
        24 => X"3388dd",
        25 => X"555577",
        26 => X"5544aa",
        27 => X"422433",
        28 => X"73172d",
        29 => X"e86a73",

        OTHERS => (OTHERS => 'U')
    );

    TYPE tile_rom_type IS ARRAY(0 TO 2 ** 13 - 1) OF unsigned(4 DOWNTO 0);
    CONSTANT tile_rom_data : tile_rom_type := (
        -- 0: grass
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011", "00011",
        OTHERS => (OTHERS => 'U')
    );

    SIGNAL palette_index : unsigned(4 DOWNTO 0); -- max 32 colors
BEGIN
    PROCESS (address)
    BEGIN
        -- get palette index from memory
        palette_index <= tile_rom_data(to_integer(address));
        data_out <= palette_rom(to_integer(palette_index));
    END PROCESS;
END ARCHITECTURE;